VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tri_144x78_2r4w
  CLASS BLOCK ;
  FOREIGN tri_144x78_2r4w ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 1500.000 ;
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.000 -0.600 4.600 3.400 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 -0.600 8.600 3.400 ;
    END
  END gnd
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.000 -0.600 12.600 3.400 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.000 -0.600 16.600 3.400 ;
    END
  END rst
  PIN delay_lclkr_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.000 -0.600 20.600 3.400 ;
    END
  END delay_lclkr_dc
  PIN mpw1_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.000 -0.600 24.600 3.400 ;
    END
  END mpw1_dc_b
  PIN mpw2_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.000 -0.600 28.600 3.400 ;
    END
  END mpw2_dc_b
  PIN func_sl_force
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.000 -0.600 32.600 3.400 ;
    END
  END func_sl_force
  PIN func_sl_thold_0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 -0.600 36.600 3.400 ;
    END
  END func_sl_thold_0_b
  PIN func_slp_sl_force
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.000 -0.600 40.600 3.400 ;
    END
  END func_slp_sl_force
  PIN func_slp_sl_thold_0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.000 -0.600 44.600 3.400 ;
    END
  END func_slp_sl_thold_0_b
  PIN sg_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.000 -0.600 48.600 3.400 ;
    END
  END sg_0
  PIN scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.000 -0.600 52.600 3.400 ;
    END
  END scan_in
  PIN scan_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 -0.600 56.600 3.400 ;
    END
  END scan_out
  PIN r_late_en_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.000 0.000 4.600 ;
    END
  END r_late_en_1
  PIN r_addr_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.000 0.000 8.600 ;
    END
  END r_addr_in_1[0]
  PIN r_addr_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.000 0.000 12.600 ;
    END
  END r_addr_in_1[1]
  PIN r_addr_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 16.000 0.000 16.600 ;
    END
  END r_addr_in_1[2]
  PIN r_addr_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 20.000 0.000 20.600 ;
    END
  END r_addr_in_1[3]
  PIN r_addr_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 24.000 0.000 24.600 ;
    END
  END r_addr_in_1[4]
  PIN r_addr_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 28.000 0.000 28.600 ;
    END
  END r_addr_in_1[5]
  PIN r_data_out_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 4.000 504.000 4.600 ;
    END
  END r_data_out_1[0]
  PIN r_data_out_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 8.000 504.000 8.600 ;
    END
  END r_data_out_1[1]
  PIN r_data_out_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 12.000 504.000 12.600 ;
    END
  END r_data_out_1[2]
  PIN r_data_out_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 16.000 504.000 16.600 ;
    END
  END r_data_out_1[3]
  PIN r_data_out_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 20.000 504.000 20.600 ;
    END
  END r_data_out_1[4]
  PIN r_data_out_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 24.000 504.000 24.600 ;
    END
  END r_data_out_1[5]
  PIN r_data_out_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 28.000 504.000 28.600 ;
    END
  END r_data_out_1[6]
  PIN r_data_out_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 32.000 504.000 32.600 ;
    END
  END r_data_out_1[7]
  PIN r_data_out_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 36.000 504.000 36.600 ;
    END
  END r_data_out_1[8]
  PIN r_data_out_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 40.000 504.000 40.600 ;
    END
  END r_data_out_1[9]
  PIN r_data_out_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 44.000 504.000 44.600 ;
    END
  END r_data_out_1[10]
  PIN r_data_out_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 48.000 504.000 48.600 ;
    END
  END r_data_out_1[11]
  PIN r_data_out_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 52.000 504.000 52.600 ;
    END
  END r_data_out_1[12]
  PIN r_data_out_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 56.000 504.000 56.600 ;
    END
  END r_data_out_1[13]
  PIN r_data_out_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 60.000 504.000 60.600 ;
    END
  END r_data_out_1[14]
  PIN r_data_out_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 64.000 504.000 64.600 ;
    END
  END r_data_out_1[15]
  PIN r_data_out_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 68.000 504.000 68.600 ;
    END
  END r_data_out_1[16]
  PIN r_data_out_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 72.000 504.000 72.600 ;
    END
  END r_data_out_1[17]
  PIN r_data_out_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 76.000 504.000 76.600 ;
    END
  END r_data_out_1[18]
  PIN r_data_out_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 80.000 504.000 80.600 ;
    END
  END r_data_out_1[19]
  PIN r_data_out_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 84.000 504.000 84.600 ;
    END
  END r_data_out_1[20]
  PIN r_data_out_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 88.000 504.000 88.600 ;
    END
  END r_data_out_1[21]
  PIN r_data_out_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 92.000 504.000 92.600 ;
    END
  END r_data_out_1[22]
  PIN r_data_out_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 96.000 504.000 96.600 ;
    END
  END r_data_out_1[23]
  PIN r_data_out_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 100.000 504.000 100.600 ;
    END
  END r_data_out_1[24]
  PIN r_data_out_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 104.000 504.000 104.600 ;
    END
  END r_data_out_1[25]
  PIN r_data_out_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 108.000 504.000 108.600 ;
    END
  END r_data_out_1[26]
  PIN r_data_out_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 112.000 504.000 112.600 ;
    END
  END r_data_out_1[27]
  PIN r_data_out_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 116.000 504.000 116.600 ;
    END
  END r_data_out_1[28]
  PIN r_data_out_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 120.000 504.000 120.600 ;
    END
  END r_data_out_1[29]
  PIN r_data_out_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 124.000 504.000 124.600 ;
    END
  END r_data_out_1[30]
  PIN r_data_out_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 128.000 504.000 128.600 ;
    END
  END r_data_out_1[31]
  PIN r_data_out_1[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 132.000 504.000 132.600 ;
    END
  END r_data_out_1[32]
  PIN r_data_out_1[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 136.000 504.000 136.600 ;
    END
  END r_data_out_1[33]
  PIN r_data_out_1[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 140.000 504.000 140.600 ;
    END
  END r_data_out_1[34]
  PIN r_data_out_1[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 144.000 504.000 144.600 ;
    END
  END r_data_out_1[35]
  PIN r_data_out_1[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 148.000 504.000 148.600 ;
    END
  END r_data_out_1[36]
  PIN r_data_out_1[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 152.000 504.000 152.600 ;
    END
  END r_data_out_1[37]
  PIN r_data_out_1[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 156.000 504.000 156.600 ;
    END
  END r_data_out_1[38]
  PIN r_data_out_1[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 160.000 504.000 160.600 ;
    END
  END r_data_out_1[39]
  PIN r_data_out_1[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 164.000 504.000 164.600 ;
    END
  END r_data_out_1[40]
  PIN r_data_out_1[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 168.000 504.000 168.600 ;
    END
  END r_data_out_1[41]
  PIN r_data_out_1[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 172.000 504.000 172.600 ;
    END
  END r_data_out_1[42]
  PIN r_data_out_1[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 176.000 504.000 176.600 ;
    END
  END r_data_out_1[43]
  PIN r_data_out_1[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 180.000 504.000 180.600 ;
    END
  END r_data_out_1[44]
  PIN r_data_out_1[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 184.000 504.000 184.600 ;
    END
  END r_data_out_1[45]
  PIN r_data_out_1[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 188.000 504.000 188.600 ;
    END
  END r_data_out_1[46]
  PIN r_data_out_1[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 192.000 504.000 192.600 ;
    END
  END r_data_out_1[47]
  PIN r_data_out_1[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 196.000 504.000 196.600 ;
    END
  END r_data_out_1[48]
  PIN r_data_out_1[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 200.000 504.000 200.600 ;
    END
  END r_data_out_1[49]
  PIN r_data_out_1[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 204.000 504.000 204.600 ;
    END
  END r_data_out_1[50]
  PIN r_data_out_1[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 208.000 504.000 208.600 ;
    END
  END r_data_out_1[51]
  PIN r_data_out_1[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 212.000 504.000 212.600 ;
    END
  END r_data_out_1[52]
  PIN r_data_out_1[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 216.000 504.000 216.600 ;
    END
  END r_data_out_1[53]
  PIN r_data_out_1[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 220.000 504.000 220.600 ;
    END
  END r_data_out_1[54]
  PIN r_data_out_1[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 224.000 504.000 224.600 ;
    END
  END r_data_out_1[55]
  PIN r_data_out_1[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 228.000 504.000 228.600 ;
    END
  END r_data_out_1[56]
  PIN r_data_out_1[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 232.000 504.000 232.600 ;
    END
  END r_data_out_1[57]
  PIN r_data_out_1[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 236.000 504.000 236.600 ;
    END
  END r_data_out_1[58]
  PIN r_data_out_1[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 240.000 504.000 240.600 ;
    END
  END r_data_out_1[59]
  PIN r_data_out_1[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 244.000 504.000 244.600 ;
    END
  END r_data_out_1[60]
  PIN r_data_out_1[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 248.000 504.000 248.600 ;
    END
  END r_data_out_1[61]
  PIN r_data_out_1[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 252.000 504.000 252.600 ;
    END
  END r_data_out_1[62]
  PIN r_data_out_1[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 256.000 504.000 256.600 ;
    END
  END r_data_out_1[63]
  PIN r_data_out_1[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 260.000 504.000 260.600 ;
    END
  END r_data_out_1[64]
  PIN r_data_out_1[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 264.000 504.000 264.600 ;
    END
  END r_data_out_1[65]
  PIN r_data_out_1[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 268.000 504.000 268.600 ;
    END
  END r_data_out_1[66]
  PIN r_data_out_1[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 272.000 504.000 272.600 ;
    END
  END r_data_out_1[67]
  PIN r_data_out_1[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 276.000 504.000 276.600 ;
    END
  END r_data_out_1[68]
  PIN r_data_out_1[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 280.000 504.000 280.600 ;
    END
  END r_data_out_1[69]
  PIN r_data_out_1[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 284.000 504.000 284.600 ;
    END
  END r_data_out_1[70]
  PIN r_data_out_1[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 288.000 504.000 288.600 ;
    END
  END r_data_out_1[71]
  PIN r_data_out_1[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 292.000 504.000 292.600 ;
    END
  END r_data_out_1[72]
  PIN r_data_out_1[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 296.000 504.000 296.600 ;
    END
  END r_data_out_1[73]
  PIN r_data_out_1[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 300.000 504.000 300.600 ;
    END
  END r_data_out_1[74]
  PIN r_data_out_1[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 304.000 504.000 304.600 ;
    END
  END r_data_out_1[75]
  PIN r_data_out_1[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 308.000 504.000 308.600 ;
    END
  END r_data_out_1[76]
  PIN r_data_out_1[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 312.000 504.000 312.600 ;
    END
  END r_data_out_1[77]
  PIN r_late_en_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 0.000 32.600 ;
    END
  END r_late_en_2
  PIN r_addr_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.000 0.000 36.600 ;
    END
  END r_addr_in_2[0]
  PIN r_addr_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.000 0.000 40.600 ;
    END
  END r_addr_in_2[1]
  PIN r_addr_in_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.000 0.000 44.600 ;
    END
  END r_addr_in_2[2]
  PIN r_addr_in_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.000 0.000 48.600 ;
    END
  END r_addr_in_2[3]
  PIN r_addr_in_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 52.000 0.000 52.600 ;
    END
  END r_addr_in_2[4]
  PIN r_addr_in_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 56.000 0.000 56.600 ;
    END
  END r_addr_in_2[5]
  PIN r_data_out_2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 316.000 504.000 316.600 ;
    END
  END r_data_out_2[0]
  PIN r_data_out_2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 320.000 504.000 320.600 ;
    END
  END r_data_out_2[1]
  PIN r_data_out_2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 324.000 504.000 324.600 ;
    END
  END r_data_out_2[2]
  PIN r_data_out_2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 328.000 504.000 328.600 ;
    END
  END r_data_out_2[3]
  PIN r_data_out_2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 332.000 504.000 332.600 ;
    END
  END r_data_out_2[4]
  PIN r_data_out_2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 336.000 504.000 336.600 ;
    END
  END r_data_out_2[5]
  PIN r_data_out_2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 340.000 504.000 340.600 ;
    END
  END r_data_out_2[6]
  PIN r_data_out_2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 344.000 504.000 344.600 ;
    END
  END r_data_out_2[7]
  PIN r_data_out_2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 348.000 504.000 348.600 ;
    END
  END r_data_out_2[8]
  PIN r_data_out_2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 352.000 504.000 352.600 ;
    END
  END r_data_out_2[9]
  PIN r_data_out_2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 356.000 504.000 356.600 ;
    END
  END r_data_out_2[10]
  PIN r_data_out_2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 360.000 504.000 360.600 ;
    END
  END r_data_out_2[11]
  PIN r_data_out_2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 364.000 504.000 364.600 ;
    END
  END r_data_out_2[12]
  PIN r_data_out_2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 368.000 504.000 368.600 ;
    END
  END r_data_out_2[13]
  PIN r_data_out_2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 372.000 504.000 372.600 ;
    END
  END r_data_out_2[14]
  PIN r_data_out_2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 376.000 504.000 376.600 ;
    END
  END r_data_out_2[15]
  PIN r_data_out_2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 380.000 504.000 380.600 ;
    END
  END r_data_out_2[16]
  PIN r_data_out_2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 384.000 504.000 384.600 ;
    END
  END r_data_out_2[17]
  PIN r_data_out_2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 388.000 504.000 388.600 ;
    END
  END r_data_out_2[18]
  PIN r_data_out_2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 392.000 504.000 392.600 ;
    END
  END r_data_out_2[19]
  PIN r_data_out_2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 396.000 504.000 396.600 ;
    END
  END r_data_out_2[20]
  PIN r_data_out_2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 400.000 504.000 400.600 ;
    END
  END r_data_out_2[21]
  PIN r_data_out_2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 404.000 504.000 404.600 ;
    END
  END r_data_out_2[22]
  PIN r_data_out_2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 408.000 504.000 408.600 ;
    END
  END r_data_out_2[23]
  PIN r_data_out_2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 412.000 504.000 412.600 ;
    END
  END r_data_out_2[24]
  PIN r_data_out_2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 416.000 504.000 416.600 ;
    END
  END r_data_out_2[25]
  PIN r_data_out_2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 420.000 504.000 420.600 ;
    END
  END r_data_out_2[26]
  PIN r_data_out_2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 424.000 504.000 424.600 ;
    END
  END r_data_out_2[27]
  PIN r_data_out_2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 428.000 504.000 428.600 ;
    END
  END r_data_out_2[28]
  PIN r_data_out_2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 432.000 504.000 432.600 ;
    END
  END r_data_out_2[29]
  PIN r_data_out_2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 436.000 504.000 436.600 ;
    END
  END r_data_out_2[30]
  PIN r_data_out_2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 440.000 504.000 440.600 ;
    END
  END r_data_out_2[31]
  PIN r_data_out_2[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 444.000 504.000 444.600 ;
    END
  END r_data_out_2[32]
  PIN r_data_out_2[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 448.000 504.000 448.600 ;
    END
  END r_data_out_2[33]
  PIN r_data_out_2[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 452.000 504.000 452.600 ;
    END
  END r_data_out_2[34]
  PIN r_data_out_2[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 456.000 504.000 456.600 ;
    END
  END r_data_out_2[35]
  PIN r_data_out_2[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 460.000 504.000 460.600 ;
    END
  END r_data_out_2[36]
  PIN r_data_out_2[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 464.000 504.000 464.600 ;
    END
  END r_data_out_2[37]
  PIN r_data_out_2[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 468.000 504.000 468.600 ;
    END
  END r_data_out_2[38]
  PIN r_data_out_2[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 472.000 504.000 472.600 ;
    END
  END r_data_out_2[39]
  PIN r_data_out_2[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 476.000 504.000 476.600 ;
    END
  END r_data_out_2[40]
  PIN r_data_out_2[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 480.000 504.000 480.600 ;
    END
  END r_data_out_2[41]
  PIN r_data_out_2[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 484.000 504.000 484.600 ;
    END
  END r_data_out_2[42]
  PIN r_data_out_2[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 488.000 504.000 488.600 ;
    END
  END r_data_out_2[43]
  PIN r_data_out_2[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 492.000 504.000 492.600 ;
    END
  END r_data_out_2[44]
  PIN r_data_out_2[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 496.000 504.000 496.600 ;
    END
  END r_data_out_2[45]
  PIN r_data_out_2[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 500.000 504.000 500.600 ;
    END
  END r_data_out_2[46]
  PIN r_data_out_2[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 504.000 504.000 504.600 ;
    END
  END r_data_out_2[47]
  PIN r_data_out_2[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 508.000 504.000 508.600 ;
    END
  END r_data_out_2[48]
  PIN r_data_out_2[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 512.000 504.000 512.600 ;
    END
  END r_data_out_2[49]
  PIN r_data_out_2[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 516.000 504.000 516.600 ;
    END
  END r_data_out_2[50]
  PIN r_data_out_2[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 520.000 504.000 520.600 ;
    END
  END r_data_out_2[51]
  PIN r_data_out_2[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 524.000 504.000 524.600 ;
    END
  END r_data_out_2[52]
  PIN r_data_out_2[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 528.000 504.000 528.600 ;
    END
  END r_data_out_2[53]
  PIN r_data_out_2[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 532.000 504.000 532.600 ;
    END
  END r_data_out_2[54]
  PIN r_data_out_2[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 536.000 504.000 536.600 ;
    END
  END r_data_out_2[55]
  PIN r_data_out_2[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 540.000 504.000 540.600 ;
    END
  END r_data_out_2[56]
  PIN r_data_out_2[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 544.000 504.000 544.600 ;
    END
  END r_data_out_2[57]
  PIN r_data_out_2[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 548.000 504.000 548.600 ;
    END
  END r_data_out_2[58]
  PIN r_data_out_2[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 552.000 504.000 552.600 ;
    END
  END r_data_out_2[59]
  PIN r_data_out_2[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 556.000 504.000 556.600 ;
    END
  END r_data_out_2[60]
  PIN r_data_out_2[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 560.000 504.000 560.600 ;
    END
  END r_data_out_2[61]
  PIN r_data_out_2[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 564.000 504.000 564.600 ;
    END
  END r_data_out_2[62]
  PIN r_data_out_2[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 568.000 504.000 568.600 ;
    END
  END r_data_out_2[63]
  PIN r_data_out_2[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 572.000 504.000 572.600 ;
    END
  END r_data_out_2[64]
  PIN r_data_out_2[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 576.000 504.000 576.600 ;
    END
  END r_data_out_2[65]
  PIN r_data_out_2[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 580.000 504.000 580.600 ;
    END
  END r_data_out_2[66]
  PIN r_data_out_2[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 584.000 504.000 584.600 ;
    END
  END r_data_out_2[67]
  PIN r_data_out_2[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 588.000 504.000 588.600 ;
    END
  END r_data_out_2[68]
  PIN r_data_out_2[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 592.000 504.000 592.600 ;
    END
  END r_data_out_2[69]
  PIN r_data_out_2[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 596.000 504.000 596.600 ;
    END
  END r_data_out_2[70]
  PIN r_data_out_2[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 600.000 504.000 600.600 ;
    END
  END r_data_out_2[71]
  PIN r_data_out_2[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 604.000 504.000 604.600 ;
    END
  END r_data_out_2[72]
  PIN r_data_out_2[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 608.000 504.000 608.600 ;
    END
  END r_data_out_2[73]
  PIN r_data_out_2[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 612.000 504.000 612.600 ;
    END
  END r_data_out_2[74]
  PIN r_data_out_2[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 616.000 504.000 616.600 ;
    END
  END r_data_out_2[75]
  PIN r_data_out_2[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 620.000 504.000 620.600 ;
    END
  END r_data_out_2[76]
  PIN r_data_out_2[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 500.000 624.000 504.000 624.600 ;
    END
  END r_data_out_2[77]
  PIN w_late_en_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 60.000 0.000 60.600 ;
    END
  END w_late_en_1
  PIN w_addr_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 64.000 0.000 64.600 ;
    END
  END w_addr_in_1[0]
  PIN w_addr_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.000 0.000 68.600 ;
    END
  END w_addr_in_1[1]
  PIN w_addr_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.000 0.000 72.600 ;
    END
  END w_addr_in_1[2]
  PIN w_addr_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.000 0.000 76.600 ;
    END
  END w_addr_in_1[3]
  PIN w_addr_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.000 0.000 80.600 ;
    END
  END w_addr_in_1[4]
  PIN w_addr_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.000 0.000 84.600 ;
    END
  END w_addr_in_1[5]
  PIN w_data_in_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.000 0.000 88.600 ;
    END
  END w_data_in_1[0]
  PIN w_data_in_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.000 0.000 92.600 ;
    END
  END w_data_in_1[1]
  PIN w_data_in_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.000 0.000 96.600 ;
    END
  END w_data_in_1[2]
  PIN w_data_in_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.000 0.000 100.600 ;
    END
  END w_data_in_1[3]
  PIN w_data_in_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.000 0.000 104.600 ;
    END
  END w_data_in_1[4]
  PIN w_data_in_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.000 0.000 108.600 ;
    END
  END w_data_in_1[5]
  PIN w_data_in_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.000 0.000 112.600 ;
    END
  END w_data_in_1[6]
  PIN w_data_in_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 116.000 0.000 116.600 ;
    END
  END w_data_in_1[7]
  PIN w_data_in_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 120.000 0.000 120.600 ;
    END
  END w_data_in_1[8]
  PIN w_data_in_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 124.000 0.000 124.600 ;
    END
  END w_data_in_1[9]
  PIN w_data_in_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 128.000 0.000 128.600 ;
    END
  END w_data_in_1[10]
  PIN w_data_in_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 132.000 0.000 132.600 ;
    END
  END w_data_in_1[11]
  PIN w_data_in_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 136.000 0.000 136.600 ;
    END
  END w_data_in_1[12]
  PIN w_data_in_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 140.000 0.000 140.600 ;
    END
  END w_data_in_1[13]
  PIN w_data_in_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 144.000 0.000 144.600 ;
    END
  END w_data_in_1[14]
  PIN w_data_in_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 148.000 0.000 148.600 ;
    END
  END w_data_in_1[15]
  PIN w_data_in_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 152.000 0.000 152.600 ;
    END
  END w_data_in_1[16]
  PIN w_data_in_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 156.000 0.000 156.600 ;
    END
  END w_data_in_1[17]
  PIN w_data_in_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 160.000 0.000 160.600 ;
    END
  END w_data_in_1[18]
  PIN w_data_in_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 164.000 0.000 164.600 ;
    END
  END w_data_in_1[19]
  PIN w_data_in_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.000 0.000 168.600 ;
    END
  END w_data_in_1[20]
  PIN w_data_in_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.000 0.000 172.600 ;
    END
  END w_data_in_1[21]
  PIN w_data_in_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.000 0.000 176.600 ;
    END
  END w_data_in_1[22]
  PIN w_data_in_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.000 0.000 180.600 ;
    END
  END w_data_in_1[23]
  PIN w_data_in_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 184.000 0.000 184.600 ;
    END
  END w_data_in_1[24]
  PIN w_data_in_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 188.000 0.000 188.600 ;
    END
  END w_data_in_1[25]
  PIN w_data_in_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 192.000 0.000 192.600 ;
    END
  END w_data_in_1[26]
  PIN w_data_in_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 196.000 0.000 196.600 ;
    END
  END w_data_in_1[27]
  PIN w_data_in_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.000 0.000 200.600 ;
    END
  END w_data_in_1[28]
  PIN w_data_in_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.000 0.000 204.600 ;
    END
  END w_data_in_1[29]
  PIN w_data_in_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.000 0.000 208.600 ;
    END
  END w_data_in_1[30]
  PIN w_data_in_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.000 0.000 212.600 ;
    END
  END w_data_in_1[31]
  PIN w_data_in_1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.000 0.000 216.600 ;
    END
  END w_data_in_1[32]
  PIN w_data_in_1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 220.000 0.000 220.600 ;
    END
  END w_data_in_1[33]
  PIN w_data_in_1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 224.000 0.000 224.600 ;
    END
  END w_data_in_1[34]
  PIN w_data_in_1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 228.000 0.000 228.600 ;
    END
  END w_data_in_1[35]
  PIN w_data_in_1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 232.000 0.000 232.600 ;
    END
  END w_data_in_1[36]
  PIN w_data_in_1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 236.000 0.000 236.600 ;
    END
  END w_data_in_1[37]
  PIN w_data_in_1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 240.000 0.000 240.600 ;
    END
  END w_data_in_1[38]
  PIN w_data_in_1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 244.000 0.000 244.600 ;
    END
  END w_data_in_1[39]
  PIN w_data_in_1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 248.000 0.000 248.600 ;
    END
  END w_data_in_1[40]
  PIN w_data_in_1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 252.000 0.000 252.600 ;
    END
  END w_data_in_1[41]
  PIN w_data_in_1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 256.000 0.000 256.600 ;
    END
  END w_data_in_1[42]
  PIN w_data_in_1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 260.000 0.000 260.600 ;
    END
  END w_data_in_1[43]
  PIN w_data_in_1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 264.000 0.000 264.600 ;
    END
  END w_data_in_1[44]
  PIN w_data_in_1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 268.000 0.000 268.600 ;
    END
  END w_data_in_1[45]
  PIN w_data_in_1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.000 0.000 272.600 ;
    END
  END w_data_in_1[46]
  PIN w_data_in_1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.000 0.000 276.600 ;
    END
  END w_data_in_1[47]
  PIN w_data_in_1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 280.000 0.000 280.600 ;
    END
  END w_data_in_1[48]
  PIN w_data_in_1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 284.000 0.000 284.600 ;
    END
  END w_data_in_1[49]
  PIN w_data_in_1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 288.000 0.000 288.600 ;
    END
  END w_data_in_1[50]
  PIN w_data_in_1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 292.000 0.000 292.600 ;
    END
  END w_data_in_1[51]
  PIN w_data_in_1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 296.000 0.000 296.600 ;
    END
  END w_data_in_1[52]
  PIN w_data_in_1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 300.000 0.000 300.600 ;
    END
  END w_data_in_1[53]
  PIN w_data_in_1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.000 0.000 304.600 ;
    END
  END w_data_in_1[54]
  PIN w_data_in_1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 308.000 0.000 308.600 ;
    END
  END w_data_in_1[55]
  PIN w_data_in_1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.000 0.000 312.600 ;
    END
  END w_data_in_1[56]
  PIN w_data_in_1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 316.000 0.000 316.600 ;
    END
  END w_data_in_1[57]
  PIN w_data_in_1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 320.000 0.000 320.600 ;
    END
  END w_data_in_1[58]
  PIN w_data_in_1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 324.000 0.000 324.600 ;
    END
  END w_data_in_1[59]
  PIN w_data_in_1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 328.000 0.000 328.600 ;
    END
  END w_data_in_1[60]
  PIN w_data_in_1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 332.000 0.000 332.600 ;
    END
  END w_data_in_1[61]
  PIN w_data_in_1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 336.000 0.000 336.600 ;
    END
  END w_data_in_1[62]
  PIN w_data_in_1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 340.000 0.000 340.600 ;
    END
  END w_data_in_1[63]
  PIN w_data_in_1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 344.000 0.000 344.600 ;
    END
  END w_data_in_1[64]
  PIN w_data_in_1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 348.000 0.000 348.600 ;
    END
  END w_data_in_1[65]
  PIN w_data_in_1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 352.000 0.000 352.600 ;
    END
  END w_data_in_1[66]
  PIN w_data_in_1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 356.000 0.000 356.600 ;
    END
  END w_data_in_1[67]
  PIN w_data_in_1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 360.000 0.000 360.600 ;
    END
  END w_data_in_1[68]
  PIN w_data_in_1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 364.000 0.000 364.600 ;
    END
  END w_data_in_1[69]
  PIN w_data_in_1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 368.000 0.000 368.600 ;
    END
  END w_data_in_1[70]
  PIN w_data_in_1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 372.000 0.000 372.600 ;
    END
  END w_data_in_1[71]
  PIN w_data_in_1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 376.000 0.000 376.600 ;
    END
  END w_data_in_1[72]
  PIN w_data_in_1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 380.000 0.000 380.600 ;
    END
  END w_data_in_1[73]
  PIN w_data_in_1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 384.000 0.000 384.600 ;
    END
  END w_data_in_1[74]
  PIN w_data_in_1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 388.000 0.000 388.600 ;
    END
  END w_data_in_1[75]
  PIN w_data_in_1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 392.000 0.000 392.600 ;
    END
  END w_data_in_1[76]
  PIN w_data_in_1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 396.000 0.000 396.600 ;
    END
  END w_data_in_1[77]
  PIN w_late_en_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 400.000 0.000 400.600 ;
    END
  END w_late_en_2
  PIN w_addr_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 404.000 0.000 404.600 ;
    END
  END w_addr_in_2[0]
  PIN w_addr_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 408.000 0.000 408.600 ;
    END
  END w_addr_in_2[1]
  PIN w_addr_in_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 412.000 0.000 412.600 ;
    END
  END w_addr_in_2[2]
  PIN w_addr_in_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 416.000 0.000 416.600 ;
    END
  END w_addr_in_2[3]
  PIN w_addr_in_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 420.000 0.000 420.600 ;
    END
  END w_addr_in_2[4]
  PIN w_addr_in_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 424.000 0.000 424.600 ;
    END
  END w_addr_in_2[5]
  PIN w_data_in_2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 428.000 0.000 428.600 ;
    END
  END w_data_in_2[0]
  PIN w_data_in_2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 432.000 0.000 432.600 ;
    END
  END w_data_in_2[1]
  PIN w_data_in_2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 436.000 0.000 436.600 ;
    END
  END w_data_in_2[2]
  PIN w_data_in_2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 440.000 0.000 440.600 ;
    END
  END w_data_in_2[3]
  PIN w_data_in_2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.000 0.000 444.600 ;
    END
  END w_data_in_2[4]
  PIN w_data_in_2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 448.000 0.000 448.600 ;
    END
  END w_data_in_2[5]
  PIN w_data_in_2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 452.000 0.000 452.600 ;
    END
  END w_data_in_2[6]
  PIN w_data_in_2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 456.000 0.000 456.600 ;
    END
  END w_data_in_2[7]
  PIN w_data_in_2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 460.000 0.000 460.600 ;
    END
  END w_data_in_2[8]
  PIN w_data_in_2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 464.000 0.000 464.600 ;
    END
  END w_data_in_2[9]
  PIN w_data_in_2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 468.000 0.000 468.600 ;
    END
  END w_data_in_2[10]
  PIN w_data_in_2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 472.000 0.000 472.600 ;
    END
  END w_data_in_2[11]
  PIN w_data_in_2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 476.000 0.000 476.600 ;
    END
  END w_data_in_2[12]
  PIN w_data_in_2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 480.000 0.000 480.600 ;
    END
  END w_data_in_2[13]
  PIN w_data_in_2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 484.000 0.000 484.600 ;
    END
  END w_data_in_2[14]
  PIN w_data_in_2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 488.000 0.000 488.600 ;
    END
  END w_data_in_2[15]
  PIN w_data_in_2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 492.000 0.000 492.600 ;
    END
  END w_data_in_2[16]
  PIN w_data_in_2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 496.000 0.000 496.600 ;
    END
  END w_data_in_2[17]
  PIN w_data_in_2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 500.000 0.000 500.600 ;
    END
  END w_data_in_2[18]
  PIN w_data_in_2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 504.000 0.000 504.600 ;
    END
  END w_data_in_2[19]
  PIN w_data_in_2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 508.000 0.000 508.600 ;
    END
  END w_data_in_2[20]
  PIN w_data_in_2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 512.000 0.000 512.600 ;
    END
  END w_data_in_2[21]
  PIN w_data_in_2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 516.000 0.000 516.600 ;
    END
  END w_data_in_2[22]
  PIN w_data_in_2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 520.000 0.000 520.600 ;
    END
  END w_data_in_2[23]
  PIN w_data_in_2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 524.000 0.000 524.600 ;
    END
  END w_data_in_2[24]
  PIN w_data_in_2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 528.000 0.000 528.600 ;
    END
  END w_data_in_2[25]
  PIN w_data_in_2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 532.000 0.000 532.600 ;
    END
  END w_data_in_2[26]
  PIN w_data_in_2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 536.000 0.000 536.600 ;
    END
  END w_data_in_2[27]
  PIN w_data_in_2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 540.000 0.000 540.600 ;
    END
  END w_data_in_2[28]
  PIN w_data_in_2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 544.000 0.000 544.600 ;
    END
  END w_data_in_2[29]
  PIN w_data_in_2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 548.000 0.000 548.600 ;
    END
  END w_data_in_2[30]
  PIN w_data_in_2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 552.000 0.000 552.600 ;
    END
  END w_data_in_2[31]
  PIN w_data_in_2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.000 0.000 556.600 ;
    END
  END w_data_in_2[32]
  PIN w_data_in_2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 560.000 0.000 560.600 ;
    END
  END w_data_in_2[33]
  PIN w_data_in_2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 564.000 0.000 564.600 ;
    END
  END w_data_in_2[34]
  PIN w_data_in_2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 568.000 0.000 568.600 ;
    END
  END w_data_in_2[35]
  PIN w_data_in_2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 572.000 0.000 572.600 ;
    END
  END w_data_in_2[36]
  PIN w_data_in_2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 576.000 0.000 576.600 ;
    END
  END w_data_in_2[37]
  PIN w_data_in_2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 580.000 0.000 580.600 ;
    END
  END w_data_in_2[38]
  PIN w_data_in_2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.000 0.000 584.600 ;
    END
  END w_data_in_2[39]
  PIN w_data_in_2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 588.000 0.000 588.600 ;
    END
  END w_data_in_2[40]
  PIN w_data_in_2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 592.000 0.000 592.600 ;
    END
  END w_data_in_2[41]
  PIN w_data_in_2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 596.000 0.000 596.600 ;
    END
  END w_data_in_2[42]
  PIN w_data_in_2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 600.000 0.000 600.600 ;
    END
  END w_data_in_2[43]
  PIN w_data_in_2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 604.000 0.000 604.600 ;
    END
  END w_data_in_2[44]
  PIN w_data_in_2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 608.000 0.000 608.600 ;
    END
  END w_data_in_2[45]
  PIN w_data_in_2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 612.000 0.000 612.600 ;
    END
  END w_data_in_2[46]
  PIN w_data_in_2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 616.000 0.000 616.600 ;
    END
  END w_data_in_2[47]
  PIN w_data_in_2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 620.000 0.000 620.600 ;
    END
  END w_data_in_2[48]
  PIN w_data_in_2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 624.000 0.000 624.600 ;
    END
  END w_data_in_2[49]
  PIN w_data_in_2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 628.000 0.000 628.600 ;
    END
  END w_data_in_2[50]
  PIN w_data_in_2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 632.000 0.000 632.600 ;
    END
  END w_data_in_2[51]
  PIN w_data_in_2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 636.000 0.000 636.600 ;
    END
  END w_data_in_2[52]
  PIN w_data_in_2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 640.000 0.000 640.600 ;
    END
  END w_data_in_2[53]
  PIN w_data_in_2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 644.000 0.000 644.600 ;
    END
  END w_data_in_2[54]
  PIN w_data_in_2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 648.000 0.000 648.600 ;
    END
  END w_data_in_2[55]
  PIN w_data_in_2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 652.000 0.000 652.600 ;
    END
  END w_data_in_2[56]
  PIN w_data_in_2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 656.000 0.000 656.600 ;
    END
  END w_data_in_2[57]
  PIN w_data_in_2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 660.000 0.000 660.600 ;
    END
  END w_data_in_2[58]
  PIN w_data_in_2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 664.000 0.000 664.600 ;
    END
  END w_data_in_2[59]
  PIN w_data_in_2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 668.000 0.000 668.600 ;
    END
  END w_data_in_2[60]
  PIN w_data_in_2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 672.000 0.000 672.600 ;
    END
  END w_data_in_2[61]
  PIN w_data_in_2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 676.000 0.000 676.600 ;
    END
  END w_data_in_2[62]
  PIN w_data_in_2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 680.000 0.000 680.600 ;
    END
  END w_data_in_2[63]
  PIN w_data_in_2[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 684.000 0.000 684.600 ;
    END
  END w_data_in_2[64]
  PIN w_data_in_2[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 688.000 0.000 688.600 ;
    END
  END w_data_in_2[65]
  PIN w_data_in_2[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 692.000 0.000 692.600 ;
    END
  END w_data_in_2[66]
  PIN w_data_in_2[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 696.000 0.000 696.600 ;
    END
  END w_data_in_2[67]
  PIN w_data_in_2[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 700.000 0.000 700.600 ;
    END
  END w_data_in_2[68]
  PIN w_data_in_2[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 704.000 0.000 704.600 ;
    END
  END w_data_in_2[69]
  PIN w_data_in_2[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 708.000 0.000 708.600 ;
    END
  END w_data_in_2[70]
  PIN w_data_in_2[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 712.000 0.000 712.600 ;
    END
  END w_data_in_2[71]
  PIN w_data_in_2[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 716.000 0.000 716.600 ;
    END
  END w_data_in_2[72]
  PIN w_data_in_2[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 720.000 0.000 720.600 ;
    END
  END w_data_in_2[73]
  PIN w_data_in_2[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 724.000 0.000 724.600 ;
    END
  END w_data_in_2[74]
  PIN w_data_in_2[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 728.000 0.000 728.600 ;
    END
  END w_data_in_2[75]
  PIN w_data_in_2[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 732.000 0.000 732.600 ;
    END
  END w_data_in_2[76]
  PIN w_data_in_2[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 736.000 0.000 736.600 ;
    END
  END w_data_in_2[77]
  PIN w_late_en_3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 740.000 0.000 740.600 ;
    END
  END w_late_en_3
  PIN w_addr_in_3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 744.000 0.000 744.600 ;
    END
  END w_addr_in_3[0]
  PIN w_addr_in_3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 748.000 0.000 748.600 ;
    END
  END w_addr_in_3[1]
  PIN w_addr_in_3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 752.000 0.000 752.600 ;
    END
  END w_addr_in_3[2]
  PIN w_addr_in_3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 756.000 0.000 756.600 ;
    END
  END w_addr_in_3[3]
  PIN w_addr_in_3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 760.000 0.000 760.600 ;
    END
  END w_addr_in_3[4]
  PIN w_addr_in_3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 764.000 0.000 764.600 ;
    END
  END w_addr_in_3[5]
  PIN w_data_in_3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 768.000 0.000 768.600 ;
    END
  END w_data_in_3[0]
  PIN w_data_in_3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 772.000 0.000 772.600 ;
    END
  END w_data_in_3[1]
  PIN w_data_in_3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 776.000 0.000 776.600 ;
    END
  END w_data_in_3[2]
  PIN w_data_in_3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 780.000 0.000 780.600 ;
    END
  END w_data_in_3[3]
  PIN w_data_in_3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 784.000 0.000 784.600 ;
    END
  END w_data_in_3[4]
  PIN w_data_in_3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 788.000 0.000 788.600 ;
    END
  END w_data_in_3[5]
  PIN w_data_in_3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 792.000 0.000 792.600 ;
    END
  END w_data_in_3[6]
  PIN w_data_in_3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 796.000 0.000 796.600 ;
    END
  END w_data_in_3[7]
  PIN w_data_in_3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 800.000 0.000 800.600 ;
    END
  END w_data_in_3[8]
  PIN w_data_in_3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 804.000 0.000 804.600 ;
    END
  END w_data_in_3[9]
  PIN w_data_in_3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 808.000 0.000 808.600 ;
    END
  END w_data_in_3[10]
  PIN w_data_in_3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 812.000 0.000 812.600 ;
    END
  END w_data_in_3[11]
  PIN w_data_in_3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 816.000 0.000 816.600 ;
    END
  END w_data_in_3[12]
  PIN w_data_in_3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 820.000 0.000 820.600 ;
    END
  END w_data_in_3[13]
  PIN w_data_in_3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 824.000 0.000 824.600 ;
    END
  END w_data_in_3[14]
  PIN w_data_in_3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 828.000 0.000 828.600 ;
    END
  END w_data_in_3[15]
  PIN w_data_in_3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 832.000 0.000 832.600 ;
    END
  END w_data_in_3[16]
  PIN w_data_in_3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 836.000 0.000 836.600 ;
    END
  END w_data_in_3[17]
  PIN w_data_in_3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 840.000 0.000 840.600 ;
    END
  END w_data_in_3[18]
  PIN w_data_in_3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 844.000 0.000 844.600 ;
    END
  END w_data_in_3[19]
  PIN w_data_in_3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 848.000 0.000 848.600 ;
    END
  END w_data_in_3[20]
  PIN w_data_in_3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 852.000 0.000 852.600 ;
    END
  END w_data_in_3[21]
  PIN w_data_in_3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 856.000 0.000 856.600 ;
    END
  END w_data_in_3[22]
  PIN w_data_in_3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 860.000 0.000 860.600 ;
    END
  END w_data_in_3[23]
  PIN w_data_in_3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 864.000 0.000 864.600 ;
    END
  END w_data_in_3[24]
  PIN w_data_in_3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 868.000 0.000 868.600 ;
    END
  END w_data_in_3[25]
  PIN w_data_in_3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 872.000 0.000 872.600 ;
    END
  END w_data_in_3[26]
  PIN w_data_in_3[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 876.000 0.000 876.600 ;
    END
  END w_data_in_3[27]
  PIN w_data_in_3[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 880.000 0.000 880.600 ;
    END
  END w_data_in_3[28]
  PIN w_data_in_3[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 884.000 0.000 884.600 ;
    END
  END w_data_in_3[29]
  PIN w_data_in_3[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 888.000 0.000 888.600 ;
    END
  END w_data_in_3[30]
  PIN w_data_in_3[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 892.000 0.000 892.600 ;
    END
  END w_data_in_3[31]
  PIN w_data_in_3[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 896.000 0.000 896.600 ;
    END
  END w_data_in_3[32]
  PIN w_data_in_3[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 900.000 0.000 900.600 ;
    END
  END w_data_in_3[33]
  PIN w_data_in_3[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 904.000 0.000 904.600 ;
    END
  END w_data_in_3[34]
  PIN w_data_in_3[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 908.000 0.000 908.600 ;
    END
  END w_data_in_3[35]
  PIN w_data_in_3[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 912.000 0.000 912.600 ;
    END
  END w_data_in_3[36]
  PIN w_data_in_3[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 916.000 0.000 916.600 ;
    END
  END w_data_in_3[37]
  PIN w_data_in_3[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 920.000 0.000 920.600 ;
    END
  END w_data_in_3[38]
  PIN w_data_in_3[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 924.000 0.000 924.600 ;
    END
  END w_data_in_3[39]
  PIN w_data_in_3[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 928.000 0.000 928.600 ;
    END
  END w_data_in_3[40]
  PIN w_data_in_3[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 932.000 0.000 932.600 ;
    END
  END w_data_in_3[41]
  PIN w_data_in_3[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 936.000 0.000 936.600 ;
    END
  END w_data_in_3[42]
  PIN w_data_in_3[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 940.000 0.000 940.600 ;
    END
  END w_data_in_3[43]
  PIN w_data_in_3[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 944.000 0.000 944.600 ;
    END
  END w_data_in_3[44]
  PIN w_data_in_3[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 948.000 0.000 948.600 ;
    END
  END w_data_in_3[45]
  PIN w_data_in_3[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 952.000 0.000 952.600 ;
    END
  END w_data_in_3[46]
  PIN w_data_in_3[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 956.000 0.000 956.600 ;
    END
  END w_data_in_3[47]
  PIN w_data_in_3[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 960.000 0.000 960.600 ;
    END
  END w_data_in_3[48]
  PIN w_data_in_3[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 964.000 0.000 964.600 ;
    END
  END w_data_in_3[49]
  PIN w_data_in_3[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 968.000 0.000 968.600 ;
    END
  END w_data_in_3[50]
  PIN w_data_in_3[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 972.000 0.000 972.600 ;
    END
  END w_data_in_3[51]
  PIN w_data_in_3[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 976.000 0.000 976.600 ;
    END
  END w_data_in_3[52]
  PIN w_data_in_3[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 980.000 0.000 980.600 ;
    END
  END w_data_in_3[53]
  PIN w_data_in_3[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 984.000 0.000 984.600 ;
    END
  END w_data_in_3[54]
  PIN w_data_in_3[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 988.000 0.000 988.600 ;
    END
  END w_data_in_3[55]
  PIN w_data_in_3[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 992.000 0.000 992.600 ;
    END
  END w_data_in_3[56]
  PIN w_data_in_3[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 996.000 0.000 996.600 ;
    END
  END w_data_in_3[57]
  PIN w_data_in_3[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1000.000 0.000 1000.600 ;
    END
  END w_data_in_3[58]
  PIN w_data_in_3[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1004.000 0.000 1004.600 ;
    END
  END w_data_in_3[59]
  PIN w_data_in_3[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1008.000 0.000 1008.600 ;
    END
  END w_data_in_3[60]
  PIN w_data_in_3[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1012.000 0.000 1012.600 ;
    END
  END w_data_in_3[61]
  PIN w_data_in_3[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1016.000 0.000 1016.600 ;
    END
  END w_data_in_3[62]
  PIN w_data_in_3[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1020.000 0.000 1020.600 ;
    END
  END w_data_in_3[63]
  PIN w_data_in_3[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1024.000 0.000 1024.600 ;
    END
  END w_data_in_3[64]
  PIN w_data_in_3[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1028.000 0.000 1028.600 ;
    END
  END w_data_in_3[65]
  PIN w_data_in_3[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1032.000 0.000 1032.600 ;
    END
  END w_data_in_3[66]
  PIN w_data_in_3[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1036.000 0.000 1036.600 ;
    END
  END w_data_in_3[67]
  PIN w_data_in_3[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1040.000 0.000 1040.600 ;
    END
  END w_data_in_3[68]
  PIN w_data_in_3[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1044.000 0.000 1044.600 ;
    END
  END w_data_in_3[69]
  PIN w_data_in_3[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1048.000 0.000 1048.600 ;
    END
  END w_data_in_3[70]
  PIN w_data_in_3[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1052.000 0.000 1052.600 ;
    END
  END w_data_in_3[71]
  PIN w_data_in_3[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1056.000 0.000 1056.600 ;
    END
  END w_data_in_3[72]
  PIN w_data_in_3[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1060.000 0.000 1060.600 ;
    END
  END w_data_in_3[73]
  PIN w_data_in_3[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1064.000 0.000 1064.600 ;
    END
  END w_data_in_3[74]
  PIN w_data_in_3[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1068.000 0.000 1068.600 ;
    END
  END w_data_in_3[75]
  PIN w_data_in_3[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1072.000 0.000 1072.600 ;
    END
  END w_data_in_3[76]
  PIN w_data_in_3[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1076.000 0.000 1076.600 ;
    END
  END w_data_in_3[77]
  PIN w_late_en_4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1080.000 0.000 1080.600 ;
    END
  END w_late_en_4
  PIN w_addr_in_4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1084.000 0.000 1084.600 ;
    END
  END w_addr_in_4[0]
  PIN w_addr_in_4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1088.000 0.000 1088.600 ;
    END
  END w_addr_in_4[1]
  PIN w_addr_in_4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1092.000 0.000 1092.600 ;
    END
  END w_addr_in_4[2]
  PIN w_addr_in_4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1096.000 0.000 1096.600 ;
    END
  END w_addr_in_4[3]
  PIN w_addr_in_4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1100.000 0.000 1100.600 ;
    END
  END w_addr_in_4[4]
  PIN w_addr_in_4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1104.000 0.000 1104.600 ;
    END
  END w_addr_in_4[5]
  PIN w_data_in_4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1108.000 0.000 1108.600 ;
    END
  END w_data_in_4[0]
  PIN w_data_in_4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1112.000 0.000 1112.600 ;
    END
  END w_data_in_4[1]
  PIN w_data_in_4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1116.000 0.000 1116.600 ;
    END
  END w_data_in_4[2]
  PIN w_data_in_4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1120.000 0.000 1120.600 ;
    END
  END w_data_in_4[3]
  PIN w_data_in_4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1124.000 0.000 1124.600 ;
    END
  END w_data_in_4[4]
  PIN w_data_in_4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1128.000 0.000 1128.600 ;
    END
  END w_data_in_4[5]
  PIN w_data_in_4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1132.000 0.000 1132.600 ;
    END
  END w_data_in_4[6]
  PIN w_data_in_4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1136.000 0.000 1136.600 ;
    END
  END w_data_in_4[7]
  PIN w_data_in_4[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1140.000 0.000 1140.600 ;
    END
  END w_data_in_4[8]
  PIN w_data_in_4[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1144.000 0.000 1144.600 ;
    END
  END w_data_in_4[9]
  PIN w_data_in_4[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1148.000 0.000 1148.600 ;
    END
  END w_data_in_4[10]
  PIN w_data_in_4[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1152.000 0.000 1152.600 ;
    END
  END w_data_in_4[11]
  PIN w_data_in_4[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1156.000 0.000 1156.600 ;
    END
  END w_data_in_4[12]
  PIN w_data_in_4[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1160.000 0.000 1160.600 ;
    END
  END w_data_in_4[13]
  PIN w_data_in_4[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1164.000 0.000 1164.600 ;
    END
  END w_data_in_4[14]
  PIN w_data_in_4[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1168.000 0.000 1168.600 ;
    END
  END w_data_in_4[15]
  PIN w_data_in_4[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1172.000 0.000 1172.600 ;
    END
  END w_data_in_4[16]
  PIN w_data_in_4[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1176.000 0.000 1176.600 ;
    END
  END w_data_in_4[17]
  PIN w_data_in_4[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1180.000 0.000 1180.600 ;
    END
  END w_data_in_4[18]
  PIN w_data_in_4[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1184.000 0.000 1184.600 ;
    END
  END w_data_in_4[19]
  PIN w_data_in_4[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1188.000 0.000 1188.600 ;
    END
  END w_data_in_4[20]
  PIN w_data_in_4[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1192.000 0.000 1192.600 ;
    END
  END w_data_in_4[21]
  PIN w_data_in_4[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1196.000 0.000 1196.600 ;
    END
  END w_data_in_4[22]
  PIN w_data_in_4[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1200.000 0.000 1200.600 ;
    END
  END w_data_in_4[23]
  PIN w_data_in_4[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1204.000 0.000 1204.600 ;
    END
  END w_data_in_4[24]
  PIN w_data_in_4[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1208.000 0.000 1208.600 ;
    END
  END w_data_in_4[25]
  PIN w_data_in_4[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1212.000 0.000 1212.600 ;
    END
  END w_data_in_4[26]
  PIN w_data_in_4[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1216.000 0.000 1216.600 ;
    END
  END w_data_in_4[27]
  PIN w_data_in_4[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1220.000 0.000 1220.600 ;
    END
  END w_data_in_4[28]
  PIN w_data_in_4[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1224.000 0.000 1224.600 ;
    END
  END w_data_in_4[29]
  PIN w_data_in_4[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1228.000 0.000 1228.600 ;
    END
  END w_data_in_4[30]
  PIN w_data_in_4[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1232.000 0.000 1232.600 ;
    END
  END w_data_in_4[31]
  PIN w_data_in_4[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1236.000 0.000 1236.600 ;
    END
  END w_data_in_4[32]
  PIN w_data_in_4[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1240.000 0.000 1240.600 ;
    END
  END w_data_in_4[33]
  PIN w_data_in_4[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1244.000 0.000 1244.600 ;
    END
  END w_data_in_4[34]
  PIN w_data_in_4[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1248.000 0.000 1248.600 ;
    END
  END w_data_in_4[35]
  PIN w_data_in_4[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1252.000 0.000 1252.600 ;
    END
  END w_data_in_4[36]
  PIN w_data_in_4[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1256.000 0.000 1256.600 ;
    END
  END w_data_in_4[37]
  PIN w_data_in_4[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1260.000 0.000 1260.600 ;
    END
  END w_data_in_4[38]
  PIN w_data_in_4[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1264.000 0.000 1264.600 ;
    END
  END w_data_in_4[39]
  PIN w_data_in_4[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1268.000 0.000 1268.600 ;
    END
  END w_data_in_4[40]
  PIN w_data_in_4[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1272.000 0.000 1272.600 ;
    END
  END w_data_in_4[41]
  PIN w_data_in_4[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1276.000 0.000 1276.600 ;
    END
  END w_data_in_4[42]
  PIN w_data_in_4[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1280.000 0.000 1280.600 ;
    END
  END w_data_in_4[43]
  PIN w_data_in_4[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1284.000 0.000 1284.600 ;
    END
  END w_data_in_4[44]
  PIN w_data_in_4[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1288.000 0.000 1288.600 ;
    END
  END w_data_in_4[45]
  PIN w_data_in_4[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1292.000 0.000 1292.600 ;
    END
  END w_data_in_4[46]
  PIN w_data_in_4[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1296.000 0.000 1296.600 ;
    END
  END w_data_in_4[47]
  PIN w_data_in_4[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1300.000 0.000 1300.600 ;
    END
  END w_data_in_4[48]
  PIN w_data_in_4[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1304.000 0.000 1304.600 ;
    END
  END w_data_in_4[49]
  PIN w_data_in_4[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1308.000 0.000 1308.600 ;
    END
  END w_data_in_4[50]
  PIN w_data_in_4[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1312.000 0.000 1312.600 ;
    END
  END w_data_in_4[51]
  PIN w_data_in_4[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1316.000 0.000 1316.600 ;
    END
  END w_data_in_4[52]
  PIN w_data_in_4[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1320.000 0.000 1320.600 ;
    END
  END w_data_in_4[53]
  PIN w_data_in_4[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1324.000 0.000 1324.600 ;
    END
  END w_data_in_4[54]
  PIN w_data_in_4[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1328.000 0.000 1328.600 ;
    END
  END w_data_in_4[55]
  PIN w_data_in_4[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1332.000 0.000 1332.600 ;
    END
  END w_data_in_4[56]
  PIN w_data_in_4[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1336.000 0.000 1336.600 ;
    END
  END w_data_in_4[57]
  PIN w_data_in_4[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1340.000 0.000 1340.600 ;
    END
  END w_data_in_4[58]
  PIN w_data_in_4[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1344.000 0.000 1344.600 ;
    END
  END w_data_in_4[59]
  PIN w_data_in_4[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1348.000 0.000 1348.600 ;
    END
  END w_data_in_4[60]
  PIN w_data_in_4[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1352.000 0.000 1352.600 ;
    END
  END w_data_in_4[61]
  PIN w_data_in_4[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1356.000 0.000 1356.600 ;
    END
  END w_data_in_4[62]
  PIN w_data_in_4[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1360.000 0.000 1360.600 ;
    END
  END w_data_in_4[63]
  PIN w_data_in_4[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1364.000 0.000 1364.600 ;
    END
  END w_data_in_4[64]
  PIN w_data_in_4[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1368.000 0.000 1368.600 ;
    END
  END w_data_in_4[65]
  PIN w_data_in_4[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1372.000 0.000 1372.600 ;
    END
  END w_data_in_4[66]
  PIN w_data_in_4[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1376.000 0.000 1376.600 ;
    END
  END w_data_in_4[67]
  PIN w_data_in_4[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1380.000 0.000 1380.600 ;
    END
  END w_data_in_4[68]
  PIN w_data_in_4[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1384.000 0.000 1384.600 ;
    END
  END w_data_in_4[69]
  PIN w_data_in_4[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1388.000 0.000 1388.600 ;
    END
  END w_data_in_4[70]
  PIN w_data_in_4[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1392.000 0.000 1392.600 ;
    END
  END w_data_in_4[71]
  PIN w_data_in_4[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1396.000 0.000 1396.600 ;
    END
  END w_data_in_4[72]
  PIN w_data_in_4[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1400.000 0.000 1400.600 ;
    END
  END w_data_in_4[73]
  PIN w_data_in_4[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1404.000 0.000 1404.600 ;
    END
  END w_data_in_4[74]
  PIN w_data_in_4[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1408.000 0.000 1408.600 ;
    END
  END w_data_in_4[75]
  PIN w_data_in_4[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1412.000 0.000 1412.600 ;
    END
  END w_data_in_4[76]
  PIN w_data_in_4[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1416.000 0.000 1416.600 ;
    END
  END w_data_in_4[77]
END tri_144x78_2r4w
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO toysram_16x12
  CLASS BLOCK ;
  FOREIGN toysram_16x12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 60.000 ;
  PIN RWL0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4.000 -0.600 4.600 3.400 ;
    END
  END RWL0[0]
  PIN RWL0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.000 -0.600 5.600 3.400 ;
    END
  END RWL0[1]
  PIN RWL0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.000 -0.600 6.600 3.400 ;
    END
  END RWL0[2]
  PIN RWL0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.000 -0.600 7.600 3.400 ;
    END
  END RWL0[3]
  PIN RWL0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.000 -0.600 8.600 3.400 ;
    END
  END RWL0[4]
  PIN RWL0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.000 -0.600 9.600 3.400 ;
    END
  END RWL0[5]
  PIN RWL0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.000 -0.600 10.600 3.400 ;
    END
  END RWL0[6]
  PIN RWL0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.000 -0.600 11.600 3.400 ;
    END
  END RWL0[7]
  PIN RWL0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.000 -0.600 12.600 3.400 ;
    END
  END RWL0[8]
  PIN RWL0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 13.000 -0.600 13.600 3.400 ;
    END
  END RWL0[9]
  PIN RWL0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.000 -0.600 14.600 3.400 ;
    END
  END RWL0[10]
  PIN RWL0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 15.000 -0.600 15.600 3.400 ;
    END
  END RWL0[11]
  PIN RWL0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.000 -0.600 16.600 3.400 ;
    END
  END RWL0[12]
  PIN RWL0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.000 -0.600 17.600 3.400 ;
    END
  END RWL0[13]
  PIN RWL0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.000 -0.600 18.600 3.400 ;
    END
  END RWL0[14]
  PIN RWL0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.000 -0.600 19.600 3.400 ;
    END
  END RWL0[15]
  PIN RWL1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.000 -0.600 20.600 3.400 ;
    END
  END RWL1[0]
  PIN RWL1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 21.000 -0.600 21.600 3.400 ;
    END
  END RWL1[1]
  PIN RWL1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.000 -0.600 22.600 3.400 ;
    END
  END RWL1[2]
  PIN RWL1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.000 -0.600 23.600 3.400 ;
    END
  END RWL1[3]
  PIN RWL1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.000 -0.600 24.600 3.400 ;
    END
  END RWL1[4]
  PIN RWL1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.000 -0.600 25.600 3.400 ;
    END
  END RWL1[5]
  PIN RWL1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 26.000 -0.600 26.600 3.400 ;
    END
  END RWL1[6]
  PIN RWL1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.000 -0.600 27.600 3.400 ;
    END
  END RWL1[7]
  PIN RWL1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.000 -0.600 28.600 3.400 ;
    END
  END RWL1[8]
  PIN RWL1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 29.000 -0.600 29.600 3.400 ;
    END
  END RWL1[9]
  PIN RWL1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.000 -0.600 30.600 3.400 ;
    END
  END RWL1[10]
  PIN RWL1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.000 -0.600 31.600 3.400 ;
    END
  END RWL1[11]
  PIN RWL1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.000 -0.600 32.600 3.400 ;
    END
  END RWL1[12]
  PIN RWL1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 33.000 -0.600 33.600 3.400 ;
    END
  END RWL1[13]
  PIN RWL1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.000 -0.600 34.600 3.400 ;
    END
  END RWL1[14]
  PIN RWL1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 35.000 -0.600 35.600 3.400 ;
    END
  END RWL1[15]
  PIN WWL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.000 -0.600 36.600 3.400 ;
    END
  END WWL[0]
  PIN WWL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 37.000 -0.600 37.600 3.400 ;
    END
  END WWL[1]
  PIN WWL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.000 -0.600 38.600 3.400 ;
    END
  END WWL[2]
  PIN WWL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 39.000 -0.600 39.600 3.400 ;
    END
  END WWL[3]
  PIN WWL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.000 -0.600 40.600 3.400 ;
    END
  END WWL[4]
  PIN WWL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 41.000 -0.600 41.600 3.400 ;
    END
  END WWL[5]
  PIN WWL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 42.000 -0.600 42.600 3.400 ;
    END
  END WWL[6]
  PIN WWL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 43.000 -0.600 43.600 3.400 ;
    END
  END WWL[7]
  PIN WWL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.000 -0.600 44.600 3.400 ;
    END
  END WWL[8]
  PIN WWL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.000 -0.600 45.600 3.400 ;
    END
  END WWL[9]
  PIN WWL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.000 -0.600 46.600 3.400 ;
    END
  END WWL[10]
  PIN WWL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 47.000 -0.600 47.600 3.400 ;
    END
  END WWL[11]
  PIN WWL[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.000 -0.600 48.600 3.400 ;
    END
  END WWL[12]
  PIN WWL[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.000 -0.600 49.600 3.400 ;
    END
  END WWL[13]
  PIN WWL[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 50.000 -0.600 50.600 3.400 ;
    END
  END WWL[14]
  PIN WWL[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.000 -0.600 51.600 3.400 ;
    END
  END WWL[15]
  PIN RBL0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 4.000 84.000 4.600 ;
    END
  END RBL0[0]
  PIN RBL0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 5.000 84.000 5.600 ;
    END
  END RBL0[1]
  PIN RBL0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 6.000 84.000 6.600 ;
    END
  END RBL0[2]
  PIN RBL0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 7.000 84.000 7.600 ;
    END
  END RBL0[3]
  PIN RBL0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 8.000 84.000 8.600 ;
    END
  END RBL0[4]
  PIN RBL0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 9.000 84.000 9.600 ;
    END
  END RBL0[5]
  PIN RBL0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 10.000 84.000 10.600 ;
    END
  END RBL0[6]
  PIN RBL0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 11.000 84.000 11.600 ;
    END
  END RBL0[7]
  PIN RBL0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 12.000 84.000 12.600 ;
    END
  END RBL0[8]
  PIN RBL0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 13.000 84.000 13.600 ;
    END
  END RBL0[9]
  PIN RBL0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 14.000 84.000 14.600 ;
    END
  END RBL0[10]
  PIN RBL0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 15.000 84.000 15.600 ;
    END
  END RBL0[11]
  PIN RBL1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 16.000 84.000 16.600 ;
    END
  END RBL1[0]
  PIN RBL1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 17.000 84.000 17.600 ;
    END
  END RBL1[1]
  PIN RBL1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 18.000 84.000 18.600 ;
    END
  END RBL1[2]
  PIN RBL1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 19.000 84.000 19.600 ;
    END
  END RBL1[3]
  PIN RBL1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 20.000 84.000 20.600 ;
    END
  END RBL1[4]
  PIN RBL1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 21.000 84.000 21.600 ;
    END
  END RBL1[5]
  PIN RBL1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 22.000 84.000 22.600 ;
    END
  END RBL1[6]
  PIN RBL1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 23.000 84.000 23.600 ;
    END
  END RBL1[7]
  PIN RBL1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 24.000 84.000 24.600 ;
    END
  END RBL1[8]
  PIN RBL1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 25.000 84.000 25.600 ;
    END
  END RBL1[9]
  PIN RBL1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 26.000 84.000 26.600 ;
    END
  END RBL1[10]
  PIN RBL1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.000 27.000 84.000 27.600 ;
    END
  END RBL1[11]
  PIN WBL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.000 -0.600 52.600 3.400 ;
    END
  END WBL[0]
  PIN WBL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 53.000 -0.600 53.600 3.400 ;
    END
  END WBL[1]
  PIN WBL[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 54.000 -0.600 54.600 3.400 ;
    END
  END WBL[2]
  PIN WBL[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.000 -0.600 55.600 3.400 ;
    END
  END WBL[3]
  PIN WBL[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 -0.600 56.600 3.400 ;
    END
  END WBL[4]
  PIN WBL[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.000 -0.600 57.600 3.400 ;
    END
  END WBL[5]
  PIN WBL[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.000 -0.600 58.600 3.400 ;
    END
  END WBL[6]
  PIN WBL[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 59.000 -0.600 59.600 3.400 ;
    END
  END WBL[7]
  PIN WBL[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.000 -0.600 60.600 3.400 ;
    END
  END WBL[8]
  PIN WBL[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 61.000 -0.600 61.600 3.400 ;
    END
  END WBL[9]
  PIN WBL[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 62.000 -0.600 62.600 3.400 ;
    END
  END WBL[10]
  PIN WBL[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 63.000 -0.600 63.600 3.400 ;
    END
  END WBL[11]
  PIN WBLb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 64.000 -0.600 64.600 3.400 ;
    END
  END WBLb[0]
  PIN WBLb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.000 -0.600 65.600 3.400 ;
    END
  END WBLb[1]
  PIN WBLb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.000 -0.600 66.600 3.400 ;
    END
  END WBLb[2]
  PIN WBLb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.000 -0.600 67.600 3.400 ;
    END
  END WBLb[3]
  PIN WBLb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.000 -0.600 68.600 3.400 ;
    END
  END WBLb[4]
  PIN WBLb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 69.000 -0.600 69.600 3.400 ;
    END
  END WBLb[5]
  PIN WBLb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.000 -0.600 70.600 3.400 ;
    END
  END WBLb[6]
  PIN WBLb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.000 -0.600 71.600 3.400 ;
    END
  END WBLb[7]
  PIN WBLb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.000 -0.600 72.600 3.400 ;
    END
  END WBLb[8]
  PIN WBLb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 73.000 -0.600 73.600 3.400 ;
    END
  END WBLb[9]
  PIN WBLb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.000 -0.600 74.600 3.400 ;
    END
  END WBLb[10]
  PIN WBLb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.000 -0.600 75.600 3.400 ;
    END
  END WBLb[11]
END toysram_16x12
END LIBRARY


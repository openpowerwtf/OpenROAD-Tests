VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tri_512x162_4w_0
  CLASS BLOCK ;
  FOREIGN tri_512x162_4w_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 3000.000 ;
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.000 0.000 4.600 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.000 0.000 8.600 ;
    END
  END vdd
  PIN vcs
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.000 0.000 12.600 ;
    END
  END vcs
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 4.000 404.000 4.600 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 8.000 404.000 8.600 ;
    END
  END rst
  PIN ccflush_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 12.000 404.000 12.600 ;
    END
  END ccflush_dc
  PIN lcb_clkoff_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 16.000 404.000 16.600 ;
    END
  END lcb_clkoff_dc_b
  PIN lcb_d_mode_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 20.000 404.000 20.600 ;
    END
  END lcb_d_mode_dc
  PIN lcb_act_dis_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 24.000 404.000 24.600 ;
    END
  END lcb_act_dis_dc
  PIN lcb_ary_nsl_thold_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 28.000 404.000 28.600 ;
    END
  END lcb_ary_nsl_thold_0
  PIN lcb_sg_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 32.000 404.000 32.600 ;
    END
  END lcb_sg_1
  PIN lcb_abst_sl_thold_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 36.000 404.000 36.600 ;
    END
  END lcb_abst_sl_thold_0
  PIN lcb_func_sl_thold_0_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 40.000 404.000 40.600 ;
    END
  END lcb_func_sl_thold_0_b
  PIN func_force
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 44.000 404.000 44.600 ;
    END
  END func_force
  PIN scan_diag_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 48.000 404.000 48.600 ;
    END
  END scan_diag_dc
  PIN scan_dis_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 52.000 404.000 52.600 ;
    END
  END scan_dis_dc_b
  PIN func_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 56.000 404.000 56.600 ;
    END
  END func_scan_in
  PIN func_scan_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 16.000 0.000 16.600 ;
    END
  END func_scan_out
  PIN abst_scan_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 60.000 404.000 60.600 ;
    END
  END abst_scan_in[0]
  PIN abst_scan_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 64.000 404.000 64.600 ;
    END
  END abst_scan_in[1]
  PIN abst_scan_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 20.000 0.000 20.600 ;
    END
  END abst_scan_out[0]
  PIN abst_scan_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 24.000 0.000 24.600 ;
    END
  END abst_scan_out[1]
  PIN lcb_delay_lclkr_np_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 68.000 404.000 68.600 ;
    END
  END lcb_delay_lclkr_np_dc
  PIN ctrl_lcb_delay_lclkr_np_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 72.000 404.000 72.600 ;
    END
  END ctrl_lcb_delay_lclkr_np_dc
  PIN dibw_lcb_delay_lclkr_np_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 76.000 404.000 76.600 ;
    END
  END dibw_lcb_delay_lclkr_np_dc
  PIN ctrl_lcb_mpw1_np_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 80.000 404.000 80.600 ;
    END
  END ctrl_lcb_mpw1_np_dc_b
  PIN dibw_lcb_mpw1_np_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 84.000 404.000 84.600 ;
    END
  END dibw_lcb_mpw1_np_dc_b
  PIN lcb_mpw1_pp_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 88.000 404.000 88.600 ;
    END
  END lcb_mpw1_pp_dc_b
  PIN lcb_mpw1_2_pp_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 92.000 404.000 92.600 ;
    END
  END lcb_mpw1_2_pp_dc_b
  PIN aodo_lcb_delay_lclkr_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 96.000 404.000 96.600 ;
    END
  END aodo_lcb_delay_lclkr_dc
  PIN aodo_lcb_mpw1_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 100.000 404.000 100.600 ;
    END
  END aodo_lcb_mpw1_dc_b
  PIN aodo_lcb_mpw2_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 104.000 404.000 104.600 ;
    END
  END aodo_lcb_mpw2_dc_b
  PIN lcb_time_sg_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 108.000 404.000 108.600 ;
    END
  END lcb_time_sg_0
  PIN lcb_time_sl_thold_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 112.000 404.000 112.600 ;
    END
  END lcb_time_sl_thold_0
  PIN time_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 116.000 404.000 116.600 ;
    END
  END time_scan_in
  PIN time_scan_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 28.000 0.000 28.600 ;
    END
  END time_scan_out
  PIN bitw_abist[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 120.000 404.000 120.600 ;
    END
  END bitw_abist[0]
  PIN bitw_abist[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 124.000 404.000 124.600 ;
    END
  END bitw_abist[1]
  PIN lcb_repr_sl_thold_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 128.000 404.000 128.600 ;
    END
  END lcb_repr_sl_thold_0
  PIN lcb_repr_sg_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 132.000 404.000 132.600 ;
    END
  END lcb_repr_sg_0
  PIN repr_scan_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 136.000 404.000 136.600 ;
    END
  END repr_scan_in
  PIN repr_scan_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 0.000 32.600 ;
    END
  END repr_scan_out
  PIN tc_lbist_ary_wrt_thru_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 140.000 404.000 140.600 ;
    END
  END tc_lbist_ary_wrt_thru_dc
  PIN abist_en_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 144.000 404.000 144.600 ;
    END
  END abist_en_1
  PIN din_abist[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 148.000 404.000 148.600 ;
    END
  END din_abist[0]
  PIN din_abist[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 152.000 404.000 152.600 ;
    END
  END din_abist[1]
  PIN din_abist[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 156.000 404.000 156.600 ;
    END
  END din_abist[2]
  PIN din_abist[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 160.000 404.000 160.600 ;
    END
  END din_abist[3]
  PIN abist_cmp_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 164.000 404.000 164.600 ;
    END
  END abist_cmp_en
  PIN abist_raw_b_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 168.000 404.000 168.600 ;
    END
  END abist_raw_b_dc
  PIN data_cmp_abist[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 172.000 404.000 172.600 ;
    END
  END data_cmp_abist[0]
  PIN data_cmp_abist[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 176.000 404.000 176.600 ;
    END
  END data_cmp_abist[1]
  PIN data_cmp_abist[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 180.000 404.000 180.600 ;
    END
  END data_cmp_abist[2]
  PIN data_cmp_abist[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 184.000 404.000 184.600 ;
    END
  END data_cmp_abist[3]
  PIN addr_abist[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 188.000 404.000 188.600 ;
    END
  END addr_abist[0]
  PIN addr_abist[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 192.000 404.000 192.600 ;
    END
  END addr_abist[1]
  PIN addr_abist[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 196.000 404.000 196.600 ;
    END
  END addr_abist[2]
  PIN addr_abist[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 200.000 404.000 200.600 ;
    END
  END addr_abist[3]
  PIN addr_abist[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 204.000 404.000 204.600 ;
    END
  END addr_abist[4]
  PIN addr_abist[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 208.000 404.000 208.600 ;
    END
  END addr_abist[5]
  PIN addr_abist[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 212.000 404.000 212.600 ;
    END
  END addr_abist[6]
  PIN addr_abist[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 216.000 404.000 216.600 ;
    END
  END addr_abist[7]
  PIN addr_abist[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 220.000 404.000 220.600 ;
    END
  END addr_abist[8]
  PIN r_wb_abist
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 224.000 404.000 224.600 ;
    END
  END r_wb_abist
  PIN write_thru_en_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 228.000 404.000 228.600 ;
    END
  END write_thru_en_dc
  PIN lcb_bolt_sl_thold_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 232.000 404.000 232.600 ;
    END
  END lcb_bolt_sl_thold_0
  PIN pc_bo_enable_2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 236.000 404.000 236.600 ;
    END
  END pc_bo_enable_2
  PIN pc_bo_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 240.000 404.000 240.600 ;
    END
  END pc_bo_reset
  PIN pc_bo_unload
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 244.000 404.000 244.600 ;
    END
  END pc_bo_unload
  PIN pc_bo_repair
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 248.000 404.000 248.600 ;
    END
  END pc_bo_repair
  PIN pc_bo_shdata
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 252.000 404.000 252.600 ;
    END
  END pc_bo_shdata
  PIN pc_bo_select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 256.000 404.000 256.600 ;
    END
  END pc_bo_select[0]
  PIN pc_bo_select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 260.000 404.000 260.600 ;
    END
  END pc_bo_select[1]
  PIN bo_pc_failout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.000 0.000 36.600 ;
    END
  END bo_pc_failout[0]
  PIN bo_pc_failout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.000 0.000 40.600 ;
    END
  END bo_pc_failout[1]
  PIN bo_pc_diagloop[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.000 0.000 44.600 ;
    END
  END bo_pc_diagloop[0]
  PIN bo_pc_diagloop[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.000 0.000 48.600 ;
    END
  END bo_pc_diagloop[1]
  PIN tri_lcb_mpw1_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 264.000 404.000 264.600 ;
    END
  END tri_lcb_mpw1_dc_b
  PIN tri_lcb_mpw2_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 268.000 404.000 268.600 ;
    END
  END tri_lcb_mpw2_dc_b
  PIN tri_lcb_delay_lclkr_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 272.000 404.000 272.600 ;
    END
  END tri_lcb_delay_lclkr_dc
  PIN tri_lcb_clkoff_dc_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 276.000 404.000 276.600 ;
    END
  END tri_lcb_clkoff_dc_b
  PIN tri_lcb_act_dis_dc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 280.000 404.000 280.600 ;
    END
  END tri_lcb_act_dis_dc
  PIN read_act[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 284.000 404.000 284.600 ;
    END
  END read_act[0]
  PIN read_act[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 288.000 404.000 288.600 ;
    END
  END read_act[1]
  PIN write_act[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 292.000 404.000 292.600 ;
    END
  END write_act[0]
  PIN write_act[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 296.000 404.000 296.600 ;
    END
  END write_act[1]
  PIN write_act[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 300.000 404.000 300.600 ;
    END
  END write_act[2]
  PIN write_act[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 304.000 404.000 304.600 ;
    END
  END write_act[3]
  PIN write_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 308.000 404.000 308.600 ;
    END
  END write_enable
  PIN write_way[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 312.000 404.000 312.600 ;
    END
  END write_way[0]
  PIN write_way[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 316.000 404.000 316.600 ;
    END
  END write_way[1]
  PIN write_way[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 320.000 404.000 320.600 ;
    END
  END write_way[2]
  PIN write_way[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 324.000 404.000 324.600 ;
    END
  END write_way[3]
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 328.000 404.000 328.600 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 332.000 404.000 332.600 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 336.000 404.000 336.600 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 340.000 404.000 340.600 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 344.000 404.000 344.600 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 348.000 404.000 348.600 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 352.000 404.000 352.600 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 356.000 404.000 356.600 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 360.000 404.000 360.600 ;
    END
  END addr[8]
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 364.000 404.000 364.600 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 368.000 404.000 368.600 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 372.000 404.000 372.600 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 376.000 404.000 376.600 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 380.000 404.000 380.600 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 384.000 404.000 384.600 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 388.000 404.000 388.600 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 392.000 404.000 392.600 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 396.000 404.000 396.600 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 400.000 404.000 400.600 ;
    END
  END data_in[9]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 404.000 404.000 404.600 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 408.000 404.000 408.600 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 412.000 404.000 412.600 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 416.000 404.000 416.600 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 420.000 404.000 420.600 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 424.000 404.000 424.600 ;
    END
  END data_in[15]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 428.000 404.000 428.600 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 432.000 404.000 432.600 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 436.000 404.000 436.600 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 440.000 404.000 440.600 ;
    END
  END data_in[19]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 444.000 404.000 444.600 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 448.000 404.000 448.600 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 452.000 404.000 452.600 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 456.000 404.000 456.600 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 460.000 404.000 460.600 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 464.000 404.000 464.600 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 468.000 404.000 468.600 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 472.000 404.000 472.600 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 476.000 404.000 476.600 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 480.000 404.000 480.600 ;
    END
  END data_in[29]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 484.000 404.000 484.600 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 488.000 404.000 488.600 ;
    END
  END data_in[31]
  PIN data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 492.000 404.000 492.600 ;
    END
  END data_in[32]
  PIN data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 496.000 404.000 496.600 ;
    END
  END data_in[33]
  PIN data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 500.000 404.000 500.600 ;
    END
  END data_in[34]
  PIN data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 504.000 404.000 504.600 ;
    END
  END data_in[35]
  PIN data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 508.000 404.000 508.600 ;
    END
  END data_in[36]
  PIN data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 512.000 404.000 512.600 ;
    END
  END data_in[37]
  PIN data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 516.000 404.000 516.600 ;
    END
  END data_in[38]
  PIN data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 520.000 404.000 520.600 ;
    END
  END data_in[39]
  PIN data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 524.000 404.000 524.600 ;
    END
  END data_in[40]
  PIN data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 528.000 404.000 528.600 ;
    END
  END data_in[41]
  PIN data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 532.000 404.000 532.600 ;
    END
  END data_in[42]
  PIN data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 536.000 404.000 536.600 ;
    END
  END data_in[43]
  PIN data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 540.000 404.000 540.600 ;
    END
  END data_in[44]
  PIN data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 544.000 404.000 544.600 ;
    END
  END data_in[45]
  PIN data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 548.000 404.000 548.600 ;
    END
  END data_in[46]
  PIN data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 552.000 404.000 552.600 ;
    END
  END data_in[47]
  PIN data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 556.000 404.000 556.600 ;
    END
  END data_in[48]
  PIN data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 560.000 404.000 560.600 ;
    END
  END data_in[49]
  PIN data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 564.000 404.000 564.600 ;
    END
  END data_in[50]
  PIN data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 568.000 404.000 568.600 ;
    END
  END data_in[51]
  PIN data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 572.000 404.000 572.600 ;
    END
  END data_in[52]
  PIN data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 576.000 404.000 576.600 ;
    END
  END data_in[53]
  PIN data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 580.000 404.000 580.600 ;
    END
  END data_in[54]
  PIN data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 584.000 404.000 584.600 ;
    END
  END data_in[55]
  PIN data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 588.000 404.000 588.600 ;
    END
  END data_in[56]
  PIN data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 592.000 404.000 592.600 ;
    END
  END data_in[57]
  PIN data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 596.000 404.000 596.600 ;
    END
  END data_in[58]
  PIN data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 600.000 404.000 600.600 ;
    END
  END data_in[59]
  PIN data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 604.000 404.000 604.600 ;
    END
  END data_in[60]
  PIN data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 608.000 404.000 608.600 ;
    END
  END data_in[61]
  PIN data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 612.000 404.000 612.600 ;
    END
  END data_in[62]
  PIN data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 616.000 404.000 616.600 ;
    END
  END data_in[63]
  PIN data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 620.000 404.000 620.600 ;
    END
  END data_in[64]
  PIN data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 624.000 404.000 624.600 ;
    END
  END data_in[65]
  PIN data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 628.000 404.000 628.600 ;
    END
  END data_in[66]
  PIN data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 632.000 404.000 632.600 ;
    END
  END data_in[67]
  PIN data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 636.000 404.000 636.600 ;
    END
  END data_in[68]
  PIN data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 640.000 404.000 640.600 ;
    END
  END data_in[69]
  PIN data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 644.000 404.000 644.600 ;
    END
  END data_in[70]
  PIN data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 648.000 404.000 648.600 ;
    END
  END data_in[71]
  PIN data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 652.000 404.000 652.600 ;
    END
  END data_in[72]
  PIN data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 656.000 404.000 656.600 ;
    END
  END data_in[73]
  PIN data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 660.000 404.000 660.600 ;
    END
  END data_in[74]
  PIN data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 664.000 404.000 664.600 ;
    END
  END data_in[75]
  PIN data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 668.000 404.000 668.600 ;
    END
  END data_in[76]
  PIN data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 672.000 404.000 672.600 ;
    END
  END data_in[77]
  PIN data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 676.000 404.000 676.600 ;
    END
  END data_in[78]
  PIN data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 680.000 404.000 680.600 ;
    END
  END data_in[79]
  PIN data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 684.000 404.000 684.600 ;
    END
  END data_in[80]
  PIN data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 688.000 404.000 688.600 ;
    END
  END data_in[81]
  PIN data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 692.000 404.000 692.600 ;
    END
  END data_in[82]
  PIN data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 696.000 404.000 696.600 ;
    END
  END data_in[83]
  PIN data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 700.000 404.000 700.600 ;
    END
  END data_in[84]
  PIN data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 704.000 404.000 704.600 ;
    END
  END data_in[85]
  PIN data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 708.000 404.000 708.600 ;
    END
  END data_in[86]
  PIN data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 712.000 404.000 712.600 ;
    END
  END data_in[87]
  PIN data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 716.000 404.000 716.600 ;
    END
  END data_in[88]
  PIN data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 720.000 404.000 720.600 ;
    END
  END data_in[89]
  PIN data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 724.000 404.000 724.600 ;
    END
  END data_in[90]
  PIN data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 728.000 404.000 728.600 ;
    END
  END data_in[91]
  PIN data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 732.000 404.000 732.600 ;
    END
  END data_in[92]
  PIN data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 736.000 404.000 736.600 ;
    END
  END data_in[93]
  PIN data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 740.000 404.000 740.600 ;
    END
  END data_in[94]
  PIN data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 744.000 404.000 744.600 ;
    END
  END data_in[95]
  PIN data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 748.000 404.000 748.600 ;
    END
  END data_in[96]
  PIN data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 752.000 404.000 752.600 ;
    END
  END data_in[97]
  PIN data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 756.000 404.000 756.600 ;
    END
  END data_in[98]
  PIN data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 760.000 404.000 760.600 ;
    END
  END data_in[99]
  PIN data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 764.000 404.000 764.600 ;
    END
  END data_in[100]
  PIN data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 768.000 404.000 768.600 ;
    END
  END data_in[101]
  PIN data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 772.000 404.000 772.600 ;
    END
  END data_in[102]
  PIN data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 776.000 404.000 776.600 ;
    END
  END data_in[103]
  PIN data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 780.000 404.000 780.600 ;
    END
  END data_in[104]
  PIN data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 784.000 404.000 784.600 ;
    END
  END data_in[105]
  PIN data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 788.000 404.000 788.600 ;
    END
  END data_in[106]
  PIN data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 792.000 404.000 792.600 ;
    END
  END data_in[107]
  PIN data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 796.000 404.000 796.600 ;
    END
  END data_in[108]
  PIN data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 800.000 404.000 800.600 ;
    END
  END data_in[109]
  PIN data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 804.000 404.000 804.600 ;
    END
  END data_in[110]
  PIN data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 808.000 404.000 808.600 ;
    END
  END data_in[111]
  PIN data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 812.000 404.000 812.600 ;
    END
  END data_in[112]
  PIN data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 816.000 404.000 816.600 ;
    END
  END data_in[113]
  PIN data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 820.000 404.000 820.600 ;
    END
  END data_in[114]
  PIN data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 824.000 404.000 824.600 ;
    END
  END data_in[115]
  PIN data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 828.000 404.000 828.600 ;
    END
  END data_in[116]
  PIN data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 832.000 404.000 832.600 ;
    END
  END data_in[117]
  PIN data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 836.000 404.000 836.600 ;
    END
  END data_in[118]
  PIN data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 840.000 404.000 840.600 ;
    END
  END data_in[119]
  PIN data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 844.000 404.000 844.600 ;
    END
  END data_in[120]
  PIN data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 848.000 404.000 848.600 ;
    END
  END data_in[121]
  PIN data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 852.000 404.000 852.600 ;
    END
  END data_in[122]
  PIN data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 856.000 404.000 856.600 ;
    END
  END data_in[123]
  PIN data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 860.000 404.000 860.600 ;
    END
  END data_in[124]
  PIN data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 864.000 404.000 864.600 ;
    END
  END data_in[125]
  PIN data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 868.000 404.000 868.600 ;
    END
  END data_in[126]
  PIN data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 872.000 404.000 872.600 ;
    END
  END data_in[127]
  PIN data_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 876.000 404.000 876.600 ;
    END
  END data_in[128]
  PIN data_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 880.000 404.000 880.600 ;
    END
  END data_in[129]
  PIN data_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 884.000 404.000 884.600 ;
    END
  END data_in[130]
  PIN data_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 888.000 404.000 888.600 ;
    END
  END data_in[131]
  PIN data_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 892.000 404.000 892.600 ;
    END
  END data_in[132]
  PIN data_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 896.000 404.000 896.600 ;
    END
  END data_in[133]
  PIN data_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 900.000 404.000 900.600 ;
    END
  END data_in[134]
  PIN data_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 904.000 404.000 904.600 ;
    END
  END data_in[135]
  PIN data_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 908.000 404.000 908.600 ;
    END
  END data_in[136]
  PIN data_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 912.000 404.000 912.600 ;
    END
  END data_in[137]
  PIN data_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 916.000 404.000 916.600 ;
    END
  END data_in[138]
  PIN data_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 920.000 404.000 920.600 ;
    END
  END data_in[139]
  PIN data_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 924.000 404.000 924.600 ;
    END
  END data_in[140]
  PIN data_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 928.000 404.000 928.600 ;
    END
  END data_in[141]
  PIN data_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 932.000 404.000 932.600 ;
    END
  END data_in[142]
  PIN data_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 936.000 404.000 936.600 ;
    END
  END data_in[143]
  PIN data_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 940.000 404.000 940.600 ;
    END
  END data_in[144]
  PIN data_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 944.000 404.000 944.600 ;
    END
  END data_in[145]
  PIN data_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 948.000 404.000 948.600 ;
    END
  END data_in[146]
  PIN data_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 952.000 404.000 952.600 ;
    END
  END data_in[147]
  PIN data_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 956.000 404.000 956.600 ;
    END
  END data_in[148]
  PIN data_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 960.000 404.000 960.600 ;
    END
  END data_in[149]
  PIN data_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 964.000 404.000 964.600 ;
    END
  END data_in[150]
  PIN data_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 968.000 404.000 968.600 ;
    END
  END data_in[151]
  PIN data_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 972.000 404.000 972.600 ;
    END
  END data_in[152]
  PIN data_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 976.000 404.000 976.600 ;
    END
  END data_in[153]
  PIN data_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 980.000 404.000 980.600 ;
    END
  END data_in[154]
  PIN data_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 984.000 404.000 984.600 ;
    END
  END data_in[155]
  PIN data_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 988.000 404.000 988.600 ;
    END
  END data_in[156]
  PIN data_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 992.000 404.000 992.600 ;
    END
  END data_in[157]
  PIN data_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 996.000 404.000 996.600 ;
    END
  END data_in[158]
  PIN data_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 1000.000 404.000 1000.600 ;
    END
  END data_in[159]
  PIN data_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 1004.000 404.000 1004.600 ;
    END
  END data_in[160]
  PIN data_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.000 1008.000 404.000 1008.600 ;
    END
  END data_in[161]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 52.000 0.000 52.600 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 56.000 0.000 56.600 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 60.000 0.000 60.600 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 64.000 0.000 64.600 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.000 0.000 68.600 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.000 0.000 72.600 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.000 0.000 76.600 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.000 0.000 80.600 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.000 0.000 84.600 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.000 0.000 88.600 ;
    END
  END data_out[9]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.000 0.000 92.600 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.000 0.000 96.600 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.000 0.000 100.600 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.000 0.000 104.600 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.000 0.000 108.600 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.000 0.000 112.600 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 116.000 0.000 116.600 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 120.000 0.000 120.600 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 124.000 0.000 124.600 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 128.000 0.000 128.600 ;
    END
  END data_out[19]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 132.000 0.000 132.600 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 136.000 0.000 136.600 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 140.000 0.000 140.600 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 144.000 0.000 144.600 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 148.000 0.000 148.600 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 152.000 0.000 152.600 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 156.000 0.000 156.600 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 160.000 0.000 160.600 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 164.000 0.000 164.600 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.000 0.000 168.600 ;
    END
  END data_out[29]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.000 0.000 172.600 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.000 0.000 176.600 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.000 0.000 180.600 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 184.000 0.000 184.600 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 188.000 0.000 188.600 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 192.000 0.000 192.600 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 196.000 0.000 196.600 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.000 0.000 200.600 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.000 0.000 204.600 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.000 0.000 208.600 ;
    END
  END data_out[39]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.000 0.000 212.600 ;
    END
  END data_out[40]
  PIN data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.000 0.000 216.600 ;
    END
  END data_out[41]
  PIN data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 220.000 0.000 220.600 ;
    END
  END data_out[42]
  PIN data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 224.000 0.000 224.600 ;
    END
  END data_out[43]
  PIN data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 228.000 0.000 228.600 ;
    END
  END data_out[44]
  PIN data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 232.000 0.000 232.600 ;
    END
  END data_out[45]
  PIN data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 236.000 0.000 236.600 ;
    END
  END data_out[46]
  PIN data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 240.000 0.000 240.600 ;
    END
  END data_out[47]
  PIN data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 244.000 0.000 244.600 ;
    END
  END data_out[48]
  PIN data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 248.000 0.000 248.600 ;
    END
  END data_out[49]
  PIN data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 252.000 0.000 252.600 ;
    END
  END data_out[50]
  PIN data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 256.000 0.000 256.600 ;
    END
  END data_out[51]
  PIN data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 260.000 0.000 260.600 ;
    END
  END data_out[52]
  PIN data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 264.000 0.000 264.600 ;
    END
  END data_out[53]
  PIN data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 268.000 0.000 268.600 ;
    END
  END data_out[54]
  PIN data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.000 0.000 272.600 ;
    END
  END data_out[55]
  PIN data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.000 0.000 276.600 ;
    END
  END data_out[56]
  PIN data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 280.000 0.000 280.600 ;
    END
  END data_out[57]
  PIN data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 284.000 0.000 284.600 ;
    END
  END data_out[58]
  PIN data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 288.000 0.000 288.600 ;
    END
  END data_out[59]
  PIN data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 292.000 0.000 292.600 ;
    END
  END data_out[60]
  PIN data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 296.000 0.000 296.600 ;
    END
  END data_out[61]
  PIN data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 300.000 0.000 300.600 ;
    END
  END data_out[62]
  PIN data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.000 0.000 304.600 ;
    END
  END data_out[63]
  PIN data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 308.000 0.000 308.600 ;
    END
  END data_out[64]
  PIN data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.000 0.000 312.600 ;
    END
  END data_out[65]
  PIN data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 316.000 0.000 316.600 ;
    END
  END data_out[66]
  PIN data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 320.000 0.000 320.600 ;
    END
  END data_out[67]
  PIN data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 324.000 0.000 324.600 ;
    END
  END data_out[68]
  PIN data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 328.000 0.000 328.600 ;
    END
  END data_out[69]
  PIN data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 332.000 0.000 332.600 ;
    END
  END data_out[70]
  PIN data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 336.000 0.000 336.600 ;
    END
  END data_out[71]
  PIN data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 340.000 0.000 340.600 ;
    END
  END data_out[72]
  PIN data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 344.000 0.000 344.600 ;
    END
  END data_out[73]
  PIN data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 348.000 0.000 348.600 ;
    END
  END data_out[74]
  PIN data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 352.000 0.000 352.600 ;
    END
  END data_out[75]
  PIN data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 356.000 0.000 356.600 ;
    END
  END data_out[76]
  PIN data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 360.000 0.000 360.600 ;
    END
  END data_out[77]
  PIN data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 364.000 0.000 364.600 ;
    END
  END data_out[78]
  PIN data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 368.000 0.000 368.600 ;
    END
  END data_out[79]
  PIN data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 372.000 0.000 372.600 ;
    END
  END data_out[80]
  PIN data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 376.000 0.000 376.600 ;
    END
  END data_out[81]
  PIN data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 380.000 0.000 380.600 ;
    END
  END data_out[82]
  PIN data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 384.000 0.000 384.600 ;
    END
  END data_out[83]
  PIN data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 388.000 0.000 388.600 ;
    END
  END data_out[84]
  PIN data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 392.000 0.000 392.600 ;
    END
  END data_out[85]
  PIN data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 396.000 0.000 396.600 ;
    END
  END data_out[86]
  PIN data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 400.000 0.000 400.600 ;
    END
  END data_out[87]
  PIN data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 404.000 0.000 404.600 ;
    END
  END data_out[88]
  PIN data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 408.000 0.000 408.600 ;
    END
  END data_out[89]
  PIN data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 412.000 0.000 412.600 ;
    END
  END data_out[90]
  PIN data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 416.000 0.000 416.600 ;
    END
  END data_out[91]
  PIN data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 420.000 0.000 420.600 ;
    END
  END data_out[92]
  PIN data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 424.000 0.000 424.600 ;
    END
  END data_out[93]
  PIN data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 428.000 0.000 428.600 ;
    END
  END data_out[94]
  PIN data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 432.000 0.000 432.600 ;
    END
  END data_out[95]
  PIN data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 436.000 0.000 436.600 ;
    END
  END data_out[96]
  PIN data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 440.000 0.000 440.600 ;
    END
  END data_out[97]
  PIN data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.000 0.000 444.600 ;
    END
  END data_out[98]
  PIN data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 448.000 0.000 448.600 ;
    END
  END data_out[99]
  PIN data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 452.000 0.000 452.600 ;
    END
  END data_out[100]
  PIN data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 456.000 0.000 456.600 ;
    END
  END data_out[101]
  PIN data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 460.000 0.000 460.600 ;
    END
  END data_out[102]
  PIN data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 464.000 0.000 464.600 ;
    END
  END data_out[103]
  PIN data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 468.000 0.000 468.600 ;
    END
  END data_out[104]
  PIN data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 472.000 0.000 472.600 ;
    END
  END data_out[105]
  PIN data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 476.000 0.000 476.600 ;
    END
  END data_out[106]
  PIN data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 480.000 0.000 480.600 ;
    END
  END data_out[107]
  PIN data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 484.000 0.000 484.600 ;
    END
  END data_out[108]
  PIN data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 488.000 0.000 488.600 ;
    END
  END data_out[109]
  PIN data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 492.000 0.000 492.600 ;
    END
  END data_out[110]
  PIN data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 496.000 0.000 496.600 ;
    END
  END data_out[111]
  PIN data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 500.000 0.000 500.600 ;
    END
  END data_out[112]
  PIN data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 504.000 0.000 504.600 ;
    END
  END data_out[113]
  PIN data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 508.000 0.000 508.600 ;
    END
  END data_out[114]
  PIN data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 512.000 0.000 512.600 ;
    END
  END data_out[115]
  PIN data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 516.000 0.000 516.600 ;
    END
  END data_out[116]
  PIN data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 520.000 0.000 520.600 ;
    END
  END data_out[117]
  PIN data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 524.000 0.000 524.600 ;
    END
  END data_out[118]
  PIN data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 528.000 0.000 528.600 ;
    END
  END data_out[119]
  PIN data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 532.000 0.000 532.600 ;
    END
  END data_out[120]
  PIN data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 536.000 0.000 536.600 ;
    END
  END data_out[121]
  PIN data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 540.000 0.000 540.600 ;
    END
  END data_out[122]
  PIN data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 544.000 0.000 544.600 ;
    END
  END data_out[123]
  PIN data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 548.000 0.000 548.600 ;
    END
  END data_out[124]
  PIN data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 552.000 0.000 552.600 ;
    END
  END data_out[125]
  PIN data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.000 0.000 556.600 ;
    END
  END data_out[126]
  PIN data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 560.000 0.000 560.600 ;
    END
  END data_out[127]
  PIN data_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 564.000 0.000 564.600 ;
    END
  END data_out[128]
  PIN data_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 568.000 0.000 568.600 ;
    END
  END data_out[129]
  PIN data_out[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 572.000 0.000 572.600 ;
    END
  END data_out[130]
  PIN data_out[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 576.000 0.000 576.600 ;
    END
  END data_out[131]
  PIN data_out[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 580.000 0.000 580.600 ;
    END
  END data_out[132]
  PIN data_out[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.000 0.000 584.600 ;
    END
  END data_out[133]
  PIN data_out[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 588.000 0.000 588.600 ;
    END
  END data_out[134]
  PIN data_out[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 592.000 0.000 592.600 ;
    END
  END data_out[135]
  PIN data_out[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 596.000 0.000 596.600 ;
    END
  END data_out[136]
  PIN data_out[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 600.000 0.000 600.600 ;
    END
  END data_out[137]
  PIN data_out[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 604.000 0.000 604.600 ;
    END
  END data_out[138]
  PIN data_out[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 608.000 0.000 608.600 ;
    END
  END data_out[139]
  PIN data_out[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 612.000 0.000 612.600 ;
    END
  END data_out[140]
  PIN data_out[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 616.000 0.000 616.600 ;
    END
  END data_out[141]
  PIN data_out[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 620.000 0.000 620.600 ;
    END
  END data_out[142]
  PIN data_out[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 624.000 0.000 624.600 ;
    END
  END data_out[143]
  PIN data_out[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 628.000 0.000 628.600 ;
    END
  END data_out[144]
  PIN data_out[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 632.000 0.000 632.600 ;
    END
  END data_out[145]
  PIN data_out[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 636.000 0.000 636.600 ;
    END
  END data_out[146]
  PIN data_out[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 640.000 0.000 640.600 ;
    END
  END data_out[147]
  PIN data_out[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 644.000 0.000 644.600 ;
    END
  END data_out[148]
  PIN data_out[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 648.000 0.000 648.600 ;
    END
  END data_out[149]
  PIN data_out[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 652.000 0.000 652.600 ;
    END
  END data_out[150]
  PIN data_out[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 656.000 0.000 656.600 ;
    END
  END data_out[151]
  PIN data_out[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 660.000 0.000 660.600 ;
    END
  END data_out[152]
  PIN data_out[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 664.000 0.000 664.600 ;
    END
  END data_out[153]
  PIN data_out[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 668.000 0.000 668.600 ;
    END
  END data_out[154]
  PIN data_out[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 672.000 0.000 672.600 ;
    END
  END data_out[155]
  PIN data_out[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 676.000 0.000 676.600 ;
    END
  END data_out[156]
  PIN data_out[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 680.000 0.000 680.600 ;
    END
  END data_out[157]
  PIN data_out[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 684.000 0.000 684.600 ;
    END
  END data_out[158]
  PIN data_out[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 688.000 0.000 688.600 ;
    END
  END data_out[159]
  PIN data_out[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 692.000 0.000 692.600 ;
    END
  END data_out[160]
  PIN data_out[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 696.000 0.000 696.600 ;
    END
  END data_out[161]
  PIN data_out[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 700.000 0.000 700.600 ;
    END
  END data_out[162]
  PIN data_out[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 704.000 0.000 704.600 ;
    END
  END data_out[163]
  PIN data_out[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 708.000 0.000 708.600 ;
    END
  END data_out[164]
  PIN data_out[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 712.000 0.000 712.600 ;
    END
  END data_out[165]
  PIN data_out[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 716.000 0.000 716.600 ;
    END
  END data_out[166]
  PIN data_out[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 720.000 0.000 720.600 ;
    END
  END data_out[167]
  PIN data_out[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 724.000 0.000 724.600 ;
    END
  END data_out[168]
  PIN data_out[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 728.000 0.000 728.600 ;
    END
  END data_out[169]
  PIN data_out[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 732.000 0.000 732.600 ;
    END
  END data_out[170]
  PIN data_out[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 736.000 0.000 736.600 ;
    END
  END data_out[171]
  PIN data_out[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 740.000 0.000 740.600 ;
    END
  END data_out[172]
  PIN data_out[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 744.000 0.000 744.600 ;
    END
  END data_out[173]
  PIN data_out[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 748.000 0.000 748.600 ;
    END
  END data_out[174]
  PIN data_out[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 752.000 0.000 752.600 ;
    END
  END data_out[175]
  PIN data_out[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 756.000 0.000 756.600 ;
    END
  END data_out[176]
  PIN data_out[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 760.000 0.000 760.600 ;
    END
  END data_out[177]
  PIN data_out[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 764.000 0.000 764.600 ;
    END
  END data_out[178]
  PIN data_out[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 768.000 0.000 768.600 ;
    END
  END data_out[179]
  PIN data_out[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 772.000 0.000 772.600 ;
    END
  END data_out[180]
  PIN data_out[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 776.000 0.000 776.600 ;
    END
  END data_out[181]
  PIN data_out[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 780.000 0.000 780.600 ;
    END
  END data_out[182]
  PIN data_out[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 784.000 0.000 784.600 ;
    END
  END data_out[183]
  PIN data_out[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 788.000 0.000 788.600 ;
    END
  END data_out[184]
  PIN data_out[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 792.000 0.000 792.600 ;
    END
  END data_out[185]
  PIN data_out[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 796.000 0.000 796.600 ;
    END
  END data_out[186]
  PIN data_out[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 800.000 0.000 800.600 ;
    END
  END data_out[187]
  PIN data_out[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 804.000 0.000 804.600 ;
    END
  END data_out[188]
  PIN data_out[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 808.000 0.000 808.600 ;
    END
  END data_out[189]
  PIN data_out[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 812.000 0.000 812.600 ;
    END
  END data_out[190]
  PIN data_out[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 816.000 0.000 816.600 ;
    END
  END data_out[191]
  PIN data_out[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 820.000 0.000 820.600 ;
    END
  END data_out[192]
  PIN data_out[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 824.000 0.000 824.600 ;
    END
  END data_out[193]
  PIN data_out[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 828.000 0.000 828.600 ;
    END
  END data_out[194]
  PIN data_out[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 832.000 0.000 832.600 ;
    END
  END data_out[195]
  PIN data_out[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 836.000 0.000 836.600 ;
    END
  END data_out[196]
  PIN data_out[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 840.000 0.000 840.600 ;
    END
  END data_out[197]
  PIN data_out[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 844.000 0.000 844.600 ;
    END
  END data_out[198]
  PIN data_out[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 848.000 0.000 848.600 ;
    END
  END data_out[199]
  PIN data_out[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 852.000 0.000 852.600 ;
    END
  END data_out[200]
  PIN data_out[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 856.000 0.000 856.600 ;
    END
  END data_out[201]
  PIN data_out[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 860.000 0.000 860.600 ;
    END
  END data_out[202]
  PIN data_out[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 864.000 0.000 864.600 ;
    END
  END data_out[203]
  PIN data_out[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 868.000 0.000 868.600 ;
    END
  END data_out[204]
  PIN data_out[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 872.000 0.000 872.600 ;
    END
  END data_out[205]
  PIN data_out[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 876.000 0.000 876.600 ;
    END
  END data_out[206]
  PIN data_out[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 880.000 0.000 880.600 ;
    END
  END data_out[207]
  PIN data_out[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 884.000 0.000 884.600 ;
    END
  END data_out[208]
  PIN data_out[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 888.000 0.000 888.600 ;
    END
  END data_out[209]
  PIN data_out[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 892.000 0.000 892.600 ;
    END
  END data_out[210]
  PIN data_out[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 896.000 0.000 896.600 ;
    END
  END data_out[211]
  PIN data_out[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 900.000 0.000 900.600 ;
    END
  END data_out[212]
  PIN data_out[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 904.000 0.000 904.600 ;
    END
  END data_out[213]
  PIN data_out[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 908.000 0.000 908.600 ;
    END
  END data_out[214]
  PIN data_out[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 912.000 0.000 912.600 ;
    END
  END data_out[215]
  PIN data_out[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 916.000 0.000 916.600 ;
    END
  END data_out[216]
  PIN data_out[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 920.000 0.000 920.600 ;
    END
  END data_out[217]
  PIN data_out[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 924.000 0.000 924.600 ;
    END
  END data_out[218]
  PIN data_out[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 928.000 0.000 928.600 ;
    END
  END data_out[219]
  PIN data_out[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 932.000 0.000 932.600 ;
    END
  END data_out[220]
  PIN data_out[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 936.000 0.000 936.600 ;
    END
  END data_out[221]
  PIN data_out[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 940.000 0.000 940.600 ;
    END
  END data_out[222]
  PIN data_out[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 944.000 0.000 944.600 ;
    END
  END data_out[223]
  PIN data_out[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 948.000 0.000 948.600 ;
    END
  END data_out[224]
  PIN data_out[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 952.000 0.000 952.600 ;
    END
  END data_out[225]
  PIN data_out[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 956.000 0.000 956.600 ;
    END
  END data_out[226]
  PIN data_out[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 960.000 0.000 960.600 ;
    END
  END data_out[227]
  PIN data_out[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 964.000 0.000 964.600 ;
    END
  END data_out[228]
  PIN data_out[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 968.000 0.000 968.600 ;
    END
  END data_out[229]
  PIN data_out[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 972.000 0.000 972.600 ;
    END
  END data_out[230]
  PIN data_out[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 976.000 0.000 976.600 ;
    END
  END data_out[231]
  PIN data_out[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 980.000 0.000 980.600 ;
    END
  END data_out[232]
  PIN data_out[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 984.000 0.000 984.600 ;
    END
  END data_out[233]
  PIN data_out[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 988.000 0.000 988.600 ;
    END
  END data_out[234]
  PIN data_out[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 992.000 0.000 992.600 ;
    END
  END data_out[235]
  PIN data_out[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 996.000 0.000 996.600 ;
    END
  END data_out[236]
  PIN data_out[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1000.000 0.000 1000.600 ;
    END
  END data_out[237]
  PIN data_out[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1004.000 0.000 1004.600 ;
    END
  END data_out[238]
  PIN data_out[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1008.000 0.000 1008.600 ;
    END
  END data_out[239]
  PIN data_out[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1012.000 0.000 1012.600 ;
    END
  END data_out[240]
  PIN data_out[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1016.000 0.000 1016.600 ;
    END
  END data_out[241]
  PIN data_out[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1020.000 0.000 1020.600 ;
    END
  END data_out[242]
  PIN data_out[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1024.000 0.000 1024.600 ;
    END
  END data_out[243]
  PIN data_out[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1028.000 0.000 1028.600 ;
    END
  END data_out[244]
  PIN data_out[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1032.000 0.000 1032.600 ;
    END
  END data_out[245]
  PIN data_out[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1036.000 0.000 1036.600 ;
    END
  END data_out[246]
  PIN data_out[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1040.000 0.000 1040.600 ;
    END
  END data_out[247]
  PIN data_out[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1044.000 0.000 1044.600 ;
    END
  END data_out[248]
  PIN data_out[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1048.000 0.000 1048.600 ;
    END
  END data_out[249]
  PIN data_out[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1052.000 0.000 1052.600 ;
    END
  END data_out[250]
  PIN data_out[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1056.000 0.000 1056.600 ;
    END
  END data_out[251]
  PIN data_out[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1060.000 0.000 1060.600 ;
    END
  END data_out[252]
  PIN data_out[253]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1064.000 0.000 1064.600 ;
    END
  END data_out[253]
  PIN data_out[254]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1068.000 0.000 1068.600 ;
    END
  END data_out[254]
  PIN data_out[255]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1072.000 0.000 1072.600 ;
    END
  END data_out[255]
  PIN data_out[256]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1076.000 0.000 1076.600 ;
    END
  END data_out[256]
  PIN data_out[257]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1080.000 0.000 1080.600 ;
    END
  END data_out[257]
  PIN data_out[258]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1084.000 0.000 1084.600 ;
    END
  END data_out[258]
  PIN data_out[259]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1088.000 0.000 1088.600 ;
    END
  END data_out[259]
  PIN data_out[260]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1092.000 0.000 1092.600 ;
    END
  END data_out[260]
  PIN data_out[261]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1096.000 0.000 1096.600 ;
    END
  END data_out[261]
  PIN data_out[262]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1100.000 0.000 1100.600 ;
    END
  END data_out[262]
  PIN data_out[263]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1104.000 0.000 1104.600 ;
    END
  END data_out[263]
  PIN data_out[264]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1108.000 0.000 1108.600 ;
    END
  END data_out[264]
  PIN data_out[265]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1112.000 0.000 1112.600 ;
    END
  END data_out[265]
  PIN data_out[266]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1116.000 0.000 1116.600 ;
    END
  END data_out[266]
  PIN data_out[267]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1120.000 0.000 1120.600 ;
    END
  END data_out[267]
  PIN data_out[268]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1124.000 0.000 1124.600 ;
    END
  END data_out[268]
  PIN data_out[269]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1128.000 0.000 1128.600 ;
    END
  END data_out[269]
  PIN data_out[270]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1132.000 0.000 1132.600 ;
    END
  END data_out[270]
  PIN data_out[271]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1136.000 0.000 1136.600 ;
    END
  END data_out[271]
  PIN data_out[272]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1140.000 0.000 1140.600 ;
    END
  END data_out[272]
  PIN data_out[273]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1144.000 0.000 1144.600 ;
    END
  END data_out[273]
  PIN data_out[274]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1148.000 0.000 1148.600 ;
    END
  END data_out[274]
  PIN data_out[275]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1152.000 0.000 1152.600 ;
    END
  END data_out[275]
  PIN data_out[276]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1156.000 0.000 1156.600 ;
    END
  END data_out[276]
  PIN data_out[277]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1160.000 0.000 1160.600 ;
    END
  END data_out[277]
  PIN data_out[278]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1164.000 0.000 1164.600 ;
    END
  END data_out[278]
  PIN data_out[279]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1168.000 0.000 1168.600 ;
    END
  END data_out[279]
  PIN data_out[280]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1172.000 0.000 1172.600 ;
    END
  END data_out[280]
  PIN data_out[281]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1176.000 0.000 1176.600 ;
    END
  END data_out[281]
  PIN data_out[282]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1180.000 0.000 1180.600 ;
    END
  END data_out[282]
  PIN data_out[283]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1184.000 0.000 1184.600 ;
    END
  END data_out[283]
  PIN data_out[284]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1188.000 0.000 1188.600 ;
    END
  END data_out[284]
  PIN data_out[285]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1192.000 0.000 1192.600 ;
    END
  END data_out[285]
  PIN data_out[286]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1196.000 0.000 1196.600 ;
    END
  END data_out[286]
  PIN data_out[287]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1200.000 0.000 1200.600 ;
    END
  END data_out[287]
  PIN data_out[288]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1204.000 0.000 1204.600 ;
    END
  END data_out[288]
  PIN data_out[289]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1208.000 0.000 1208.600 ;
    END
  END data_out[289]
  PIN data_out[290]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1212.000 0.000 1212.600 ;
    END
  END data_out[290]
  PIN data_out[291]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1216.000 0.000 1216.600 ;
    END
  END data_out[291]
  PIN data_out[292]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1220.000 0.000 1220.600 ;
    END
  END data_out[292]
  PIN data_out[293]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1224.000 0.000 1224.600 ;
    END
  END data_out[293]
  PIN data_out[294]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1228.000 0.000 1228.600 ;
    END
  END data_out[294]
  PIN data_out[295]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1232.000 0.000 1232.600 ;
    END
  END data_out[295]
  PIN data_out[296]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1236.000 0.000 1236.600 ;
    END
  END data_out[296]
  PIN data_out[297]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1240.000 0.000 1240.600 ;
    END
  END data_out[297]
  PIN data_out[298]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1244.000 0.000 1244.600 ;
    END
  END data_out[298]
  PIN data_out[299]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1248.000 0.000 1248.600 ;
    END
  END data_out[299]
  PIN data_out[300]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1252.000 0.000 1252.600 ;
    END
  END data_out[300]
  PIN data_out[301]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1256.000 0.000 1256.600 ;
    END
  END data_out[301]
  PIN data_out[302]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1260.000 0.000 1260.600 ;
    END
  END data_out[302]
  PIN data_out[303]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1264.000 0.000 1264.600 ;
    END
  END data_out[303]
  PIN data_out[304]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1268.000 0.000 1268.600 ;
    END
  END data_out[304]
  PIN data_out[305]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1272.000 0.000 1272.600 ;
    END
  END data_out[305]
  PIN data_out[306]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1276.000 0.000 1276.600 ;
    END
  END data_out[306]
  PIN data_out[307]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1280.000 0.000 1280.600 ;
    END
  END data_out[307]
  PIN data_out[308]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1284.000 0.000 1284.600 ;
    END
  END data_out[308]
  PIN data_out[309]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1288.000 0.000 1288.600 ;
    END
  END data_out[309]
  PIN data_out[310]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1292.000 0.000 1292.600 ;
    END
  END data_out[310]
  PIN data_out[311]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1296.000 0.000 1296.600 ;
    END
  END data_out[311]
  PIN data_out[312]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1300.000 0.000 1300.600 ;
    END
  END data_out[312]
  PIN data_out[313]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1304.000 0.000 1304.600 ;
    END
  END data_out[313]
  PIN data_out[314]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1308.000 0.000 1308.600 ;
    END
  END data_out[314]
  PIN data_out[315]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1312.000 0.000 1312.600 ;
    END
  END data_out[315]
  PIN data_out[316]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1316.000 0.000 1316.600 ;
    END
  END data_out[316]
  PIN data_out[317]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1320.000 0.000 1320.600 ;
    END
  END data_out[317]
  PIN data_out[318]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1324.000 0.000 1324.600 ;
    END
  END data_out[318]
  PIN data_out[319]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1328.000 0.000 1328.600 ;
    END
  END data_out[319]
  PIN data_out[320]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1332.000 0.000 1332.600 ;
    END
  END data_out[320]
  PIN data_out[321]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1336.000 0.000 1336.600 ;
    END
  END data_out[321]
  PIN data_out[322]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1340.000 0.000 1340.600 ;
    END
  END data_out[322]
  PIN data_out[323]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1344.000 0.000 1344.600 ;
    END
  END data_out[323]
  PIN data_out[324]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1348.000 0.000 1348.600 ;
    END
  END data_out[324]
  PIN data_out[325]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1352.000 0.000 1352.600 ;
    END
  END data_out[325]
  PIN data_out[326]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1356.000 0.000 1356.600 ;
    END
  END data_out[326]
  PIN data_out[327]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1360.000 0.000 1360.600 ;
    END
  END data_out[327]
  PIN data_out[328]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1364.000 0.000 1364.600 ;
    END
  END data_out[328]
  PIN data_out[329]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1368.000 0.000 1368.600 ;
    END
  END data_out[329]
  PIN data_out[330]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1372.000 0.000 1372.600 ;
    END
  END data_out[330]
  PIN data_out[331]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1376.000 0.000 1376.600 ;
    END
  END data_out[331]
  PIN data_out[332]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1380.000 0.000 1380.600 ;
    END
  END data_out[332]
  PIN data_out[333]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1384.000 0.000 1384.600 ;
    END
  END data_out[333]
  PIN data_out[334]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1388.000 0.000 1388.600 ;
    END
  END data_out[334]
  PIN data_out[335]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1392.000 0.000 1392.600 ;
    END
  END data_out[335]
  PIN data_out[336]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1396.000 0.000 1396.600 ;
    END
  END data_out[336]
  PIN data_out[337]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1400.000 0.000 1400.600 ;
    END
  END data_out[337]
  PIN data_out[338]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1404.000 0.000 1404.600 ;
    END
  END data_out[338]
  PIN data_out[339]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1408.000 0.000 1408.600 ;
    END
  END data_out[339]
  PIN data_out[340]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1412.000 0.000 1412.600 ;
    END
  END data_out[340]
  PIN data_out[341]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1416.000 0.000 1416.600 ;
    END
  END data_out[341]
  PIN data_out[342]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1420.000 0.000 1420.600 ;
    END
  END data_out[342]
  PIN data_out[343]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1424.000 0.000 1424.600 ;
    END
  END data_out[343]
  PIN data_out[344]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1428.000 0.000 1428.600 ;
    END
  END data_out[344]
  PIN data_out[345]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1432.000 0.000 1432.600 ;
    END
  END data_out[345]
  PIN data_out[346]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1436.000 0.000 1436.600 ;
    END
  END data_out[346]
  PIN data_out[347]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1440.000 0.000 1440.600 ;
    END
  END data_out[347]
  PIN data_out[348]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1444.000 0.000 1444.600 ;
    END
  END data_out[348]
  PIN data_out[349]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1448.000 0.000 1448.600 ;
    END
  END data_out[349]
  PIN data_out[350]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1452.000 0.000 1452.600 ;
    END
  END data_out[350]
  PIN data_out[351]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1456.000 0.000 1456.600 ;
    END
  END data_out[351]
  PIN data_out[352]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1460.000 0.000 1460.600 ;
    END
  END data_out[352]
  PIN data_out[353]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1464.000 0.000 1464.600 ;
    END
  END data_out[353]
  PIN data_out[354]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1468.000 0.000 1468.600 ;
    END
  END data_out[354]
  PIN data_out[355]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1472.000 0.000 1472.600 ;
    END
  END data_out[355]
  PIN data_out[356]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1476.000 0.000 1476.600 ;
    END
  END data_out[356]
  PIN data_out[357]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1480.000 0.000 1480.600 ;
    END
  END data_out[357]
  PIN data_out[358]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1484.000 0.000 1484.600 ;
    END
  END data_out[358]
  PIN data_out[359]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1488.000 0.000 1488.600 ;
    END
  END data_out[359]
  PIN data_out[360]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1492.000 0.000 1492.600 ;
    END
  END data_out[360]
  PIN data_out[361]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1496.000 0.000 1496.600 ;
    END
  END data_out[361]
  PIN data_out[362]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1500.000 0.000 1500.600 ;
    END
  END data_out[362]
  PIN data_out[363]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1504.000 0.000 1504.600 ;
    END
  END data_out[363]
  PIN data_out[364]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1508.000 0.000 1508.600 ;
    END
  END data_out[364]
  PIN data_out[365]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1512.000 0.000 1512.600 ;
    END
  END data_out[365]
  PIN data_out[366]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1516.000 0.000 1516.600 ;
    END
  END data_out[366]
  PIN data_out[367]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1520.000 0.000 1520.600 ;
    END
  END data_out[367]
  PIN data_out[368]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1524.000 0.000 1524.600 ;
    END
  END data_out[368]
  PIN data_out[369]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1528.000 0.000 1528.600 ;
    END
  END data_out[369]
  PIN data_out[370]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1532.000 0.000 1532.600 ;
    END
  END data_out[370]
  PIN data_out[371]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1536.000 0.000 1536.600 ;
    END
  END data_out[371]
  PIN data_out[372]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1540.000 0.000 1540.600 ;
    END
  END data_out[372]
  PIN data_out[373]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1544.000 0.000 1544.600 ;
    END
  END data_out[373]
  PIN data_out[374]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1548.000 0.000 1548.600 ;
    END
  END data_out[374]
  PIN data_out[375]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1552.000 0.000 1552.600 ;
    END
  END data_out[375]
  PIN data_out[376]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1556.000 0.000 1556.600 ;
    END
  END data_out[376]
  PIN data_out[377]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1560.000 0.000 1560.600 ;
    END
  END data_out[377]
  PIN data_out[378]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1564.000 0.000 1564.600 ;
    END
  END data_out[378]
  PIN data_out[379]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1568.000 0.000 1568.600 ;
    END
  END data_out[379]
  PIN data_out[380]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1572.000 0.000 1572.600 ;
    END
  END data_out[380]
  PIN data_out[381]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1576.000 0.000 1576.600 ;
    END
  END data_out[381]
  PIN data_out[382]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1580.000 0.000 1580.600 ;
    END
  END data_out[382]
  PIN data_out[383]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1584.000 0.000 1584.600 ;
    END
  END data_out[383]
  PIN data_out[384]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1588.000 0.000 1588.600 ;
    END
  END data_out[384]
  PIN data_out[385]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1592.000 0.000 1592.600 ;
    END
  END data_out[385]
  PIN data_out[386]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1596.000 0.000 1596.600 ;
    END
  END data_out[386]
  PIN data_out[387]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1600.000 0.000 1600.600 ;
    END
  END data_out[387]
  PIN data_out[388]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1604.000 0.000 1604.600 ;
    END
  END data_out[388]
  PIN data_out[389]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1608.000 0.000 1608.600 ;
    END
  END data_out[389]
  PIN data_out[390]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1612.000 0.000 1612.600 ;
    END
  END data_out[390]
  PIN data_out[391]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1616.000 0.000 1616.600 ;
    END
  END data_out[391]
  PIN data_out[392]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1620.000 0.000 1620.600 ;
    END
  END data_out[392]
  PIN data_out[393]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1624.000 0.000 1624.600 ;
    END
  END data_out[393]
  PIN data_out[394]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1628.000 0.000 1628.600 ;
    END
  END data_out[394]
  PIN data_out[395]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1632.000 0.000 1632.600 ;
    END
  END data_out[395]
  PIN data_out[396]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1636.000 0.000 1636.600 ;
    END
  END data_out[396]
  PIN data_out[397]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1640.000 0.000 1640.600 ;
    END
  END data_out[397]
  PIN data_out[398]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1644.000 0.000 1644.600 ;
    END
  END data_out[398]
  PIN data_out[399]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1648.000 0.000 1648.600 ;
    END
  END data_out[399]
  PIN data_out[400]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1652.000 0.000 1652.600 ;
    END
  END data_out[400]
  PIN data_out[401]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1656.000 0.000 1656.600 ;
    END
  END data_out[401]
  PIN data_out[402]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1660.000 0.000 1660.600 ;
    END
  END data_out[402]
  PIN data_out[403]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1664.000 0.000 1664.600 ;
    END
  END data_out[403]
  PIN data_out[404]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1668.000 0.000 1668.600 ;
    END
  END data_out[404]
  PIN data_out[405]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1672.000 0.000 1672.600 ;
    END
  END data_out[405]
  PIN data_out[406]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1676.000 0.000 1676.600 ;
    END
  END data_out[406]
  PIN data_out[407]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1680.000 0.000 1680.600 ;
    END
  END data_out[407]
  PIN data_out[408]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1684.000 0.000 1684.600 ;
    END
  END data_out[408]
  PIN data_out[409]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1688.000 0.000 1688.600 ;
    END
  END data_out[409]
  PIN data_out[410]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1692.000 0.000 1692.600 ;
    END
  END data_out[410]
  PIN data_out[411]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1696.000 0.000 1696.600 ;
    END
  END data_out[411]
  PIN data_out[412]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1700.000 0.000 1700.600 ;
    END
  END data_out[412]
  PIN data_out[413]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1704.000 0.000 1704.600 ;
    END
  END data_out[413]
  PIN data_out[414]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1708.000 0.000 1708.600 ;
    END
  END data_out[414]
  PIN data_out[415]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1712.000 0.000 1712.600 ;
    END
  END data_out[415]
  PIN data_out[416]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1716.000 0.000 1716.600 ;
    END
  END data_out[416]
  PIN data_out[417]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1720.000 0.000 1720.600 ;
    END
  END data_out[417]
  PIN data_out[418]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1724.000 0.000 1724.600 ;
    END
  END data_out[418]
  PIN data_out[419]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1728.000 0.000 1728.600 ;
    END
  END data_out[419]
  PIN data_out[420]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1732.000 0.000 1732.600 ;
    END
  END data_out[420]
  PIN data_out[421]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1736.000 0.000 1736.600 ;
    END
  END data_out[421]
  PIN data_out[422]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1740.000 0.000 1740.600 ;
    END
  END data_out[422]
  PIN data_out[423]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1744.000 0.000 1744.600 ;
    END
  END data_out[423]
  PIN data_out[424]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1748.000 0.000 1748.600 ;
    END
  END data_out[424]
  PIN data_out[425]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1752.000 0.000 1752.600 ;
    END
  END data_out[425]
  PIN data_out[426]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1756.000 0.000 1756.600 ;
    END
  END data_out[426]
  PIN data_out[427]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1760.000 0.000 1760.600 ;
    END
  END data_out[427]
  PIN data_out[428]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1764.000 0.000 1764.600 ;
    END
  END data_out[428]
  PIN data_out[429]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1768.000 0.000 1768.600 ;
    END
  END data_out[429]
  PIN data_out[430]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1772.000 0.000 1772.600 ;
    END
  END data_out[430]
  PIN data_out[431]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1776.000 0.000 1776.600 ;
    END
  END data_out[431]
  PIN data_out[432]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1780.000 0.000 1780.600 ;
    END
  END data_out[432]
  PIN data_out[433]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1784.000 0.000 1784.600 ;
    END
  END data_out[433]
  PIN data_out[434]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1788.000 0.000 1788.600 ;
    END
  END data_out[434]
  PIN data_out[435]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1792.000 0.000 1792.600 ;
    END
  END data_out[435]
  PIN data_out[436]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1796.000 0.000 1796.600 ;
    END
  END data_out[436]
  PIN data_out[437]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1800.000 0.000 1800.600 ;
    END
  END data_out[437]
  PIN data_out[438]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1804.000 0.000 1804.600 ;
    END
  END data_out[438]
  PIN data_out[439]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1808.000 0.000 1808.600 ;
    END
  END data_out[439]
  PIN data_out[440]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1812.000 0.000 1812.600 ;
    END
  END data_out[440]
  PIN data_out[441]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1816.000 0.000 1816.600 ;
    END
  END data_out[441]
  PIN data_out[442]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1820.000 0.000 1820.600 ;
    END
  END data_out[442]
  PIN data_out[443]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1824.000 0.000 1824.600 ;
    END
  END data_out[443]
  PIN data_out[444]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1828.000 0.000 1828.600 ;
    END
  END data_out[444]
  PIN data_out[445]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1832.000 0.000 1832.600 ;
    END
  END data_out[445]
  PIN data_out[446]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1836.000 0.000 1836.600 ;
    END
  END data_out[446]
  PIN data_out[447]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1840.000 0.000 1840.600 ;
    END
  END data_out[447]
  PIN data_out[448]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1844.000 0.000 1844.600 ;
    END
  END data_out[448]
  PIN data_out[449]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1848.000 0.000 1848.600 ;
    END
  END data_out[449]
  PIN data_out[450]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1852.000 0.000 1852.600 ;
    END
  END data_out[450]
  PIN data_out[451]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1856.000 0.000 1856.600 ;
    END
  END data_out[451]
  PIN data_out[452]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1860.000 0.000 1860.600 ;
    END
  END data_out[452]
  PIN data_out[453]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1864.000 0.000 1864.600 ;
    END
  END data_out[453]
  PIN data_out[454]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1868.000 0.000 1868.600 ;
    END
  END data_out[454]
  PIN data_out[455]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1872.000 0.000 1872.600 ;
    END
  END data_out[455]
  PIN data_out[456]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1876.000 0.000 1876.600 ;
    END
  END data_out[456]
  PIN data_out[457]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1880.000 0.000 1880.600 ;
    END
  END data_out[457]
  PIN data_out[458]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1884.000 0.000 1884.600 ;
    END
  END data_out[458]
  PIN data_out[459]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1888.000 0.000 1888.600 ;
    END
  END data_out[459]
  PIN data_out[460]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1892.000 0.000 1892.600 ;
    END
  END data_out[460]
  PIN data_out[461]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1896.000 0.000 1896.600 ;
    END
  END data_out[461]
  PIN data_out[462]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1900.000 0.000 1900.600 ;
    END
  END data_out[462]
  PIN data_out[463]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1904.000 0.000 1904.600 ;
    END
  END data_out[463]
  PIN data_out[464]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1908.000 0.000 1908.600 ;
    END
  END data_out[464]
  PIN data_out[465]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1912.000 0.000 1912.600 ;
    END
  END data_out[465]
  PIN data_out[466]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1916.000 0.000 1916.600 ;
    END
  END data_out[466]
  PIN data_out[467]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1920.000 0.000 1920.600 ;
    END
  END data_out[467]
  PIN data_out[468]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1924.000 0.000 1924.600 ;
    END
  END data_out[468]
  PIN data_out[469]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1928.000 0.000 1928.600 ;
    END
  END data_out[469]
  PIN data_out[470]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1932.000 0.000 1932.600 ;
    END
  END data_out[470]
  PIN data_out[471]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1936.000 0.000 1936.600 ;
    END
  END data_out[471]
  PIN data_out[472]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1940.000 0.000 1940.600 ;
    END
  END data_out[472]
  PIN data_out[473]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1944.000 0.000 1944.600 ;
    END
  END data_out[473]
  PIN data_out[474]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1948.000 0.000 1948.600 ;
    END
  END data_out[474]
  PIN data_out[475]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1952.000 0.000 1952.600 ;
    END
  END data_out[475]
  PIN data_out[476]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1956.000 0.000 1956.600 ;
    END
  END data_out[476]
  PIN data_out[477]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1960.000 0.000 1960.600 ;
    END
  END data_out[477]
  PIN data_out[478]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1964.000 0.000 1964.600 ;
    END
  END data_out[478]
  PIN data_out[479]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1968.000 0.000 1968.600 ;
    END
  END data_out[479]
  PIN data_out[480]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1972.000 0.000 1972.600 ;
    END
  END data_out[480]
  PIN data_out[481]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1976.000 0.000 1976.600 ;
    END
  END data_out[481]
  PIN data_out[482]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1980.000 0.000 1980.600 ;
    END
  END data_out[482]
  PIN data_out[483]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1984.000 0.000 1984.600 ;
    END
  END data_out[483]
  PIN data_out[484]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1988.000 0.000 1988.600 ;
    END
  END data_out[484]
  PIN data_out[485]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1992.000 0.000 1992.600 ;
    END
  END data_out[485]
  PIN data_out[486]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 1996.000 0.000 1996.600 ;
    END
  END data_out[486]
  PIN data_out[487]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2000.000 0.000 2000.600 ;
    END
  END data_out[487]
  PIN data_out[488]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2004.000 0.000 2004.600 ;
    END
  END data_out[488]
  PIN data_out[489]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2008.000 0.000 2008.600 ;
    END
  END data_out[489]
  PIN data_out[490]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2012.000 0.000 2012.600 ;
    END
  END data_out[490]
  PIN data_out[491]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2016.000 0.000 2016.600 ;
    END
  END data_out[491]
  PIN data_out[492]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2020.000 0.000 2020.600 ;
    END
  END data_out[492]
  PIN data_out[493]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2024.000 0.000 2024.600 ;
    END
  END data_out[493]
  PIN data_out[494]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2028.000 0.000 2028.600 ;
    END
  END data_out[494]
  PIN data_out[495]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2032.000 0.000 2032.600 ;
    END
  END data_out[495]
  PIN data_out[496]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2036.000 0.000 2036.600 ;
    END
  END data_out[496]
  PIN data_out[497]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2040.000 0.000 2040.600 ;
    END
  END data_out[497]
  PIN data_out[498]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2044.000 0.000 2044.600 ;
    END
  END data_out[498]
  PIN data_out[499]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2048.000 0.000 2048.600 ;
    END
  END data_out[499]
  PIN data_out[500]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2052.000 0.000 2052.600 ;
    END
  END data_out[500]
  PIN data_out[501]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2056.000 0.000 2056.600 ;
    END
  END data_out[501]
  PIN data_out[502]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2060.000 0.000 2060.600 ;
    END
  END data_out[502]
  PIN data_out[503]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2064.000 0.000 2064.600 ;
    END
  END data_out[503]
  PIN data_out[504]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2068.000 0.000 2068.600 ;
    END
  END data_out[504]
  PIN data_out[505]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2072.000 0.000 2072.600 ;
    END
  END data_out[505]
  PIN data_out[506]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2076.000 0.000 2076.600 ;
    END
  END data_out[506]
  PIN data_out[507]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2080.000 0.000 2080.600 ;
    END
  END data_out[507]
  PIN data_out[508]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2084.000 0.000 2084.600 ;
    END
  END data_out[508]
  PIN data_out[509]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2088.000 0.000 2088.600 ;
    END
  END data_out[509]
  PIN data_out[510]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2092.000 0.000 2092.600 ;
    END
  END data_out[510]
  PIN data_out[511]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2096.000 0.000 2096.600 ;
    END
  END data_out[511]
  PIN data_out[512]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2100.000 0.000 2100.600 ;
    END
  END data_out[512]
  PIN data_out[513]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2104.000 0.000 2104.600 ;
    END
  END data_out[513]
  PIN data_out[514]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2108.000 0.000 2108.600 ;
    END
  END data_out[514]
  PIN data_out[515]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2112.000 0.000 2112.600 ;
    END
  END data_out[515]
  PIN data_out[516]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2116.000 0.000 2116.600 ;
    END
  END data_out[516]
  PIN data_out[517]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2120.000 0.000 2120.600 ;
    END
  END data_out[517]
  PIN data_out[518]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2124.000 0.000 2124.600 ;
    END
  END data_out[518]
  PIN data_out[519]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2128.000 0.000 2128.600 ;
    END
  END data_out[519]
  PIN data_out[520]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2132.000 0.000 2132.600 ;
    END
  END data_out[520]
  PIN data_out[521]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2136.000 0.000 2136.600 ;
    END
  END data_out[521]
  PIN data_out[522]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2140.000 0.000 2140.600 ;
    END
  END data_out[522]
  PIN data_out[523]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2144.000 0.000 2144.600 ;
    END
  END data_out[523]
  PIN data_out[524]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2148.000 0.000 2148.600 ;
    END
  END data_out[524]
  PIN data_out[525]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2152.000 0.000 2152.600 ;
    END
  END data_out[525]
  PIN data_out[526]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2156.000 0.000 2156.600 ;
    END
  END data_out[526]
  PIN data_out[527]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2160.000 0.000 2160.600 ;
    END
  END data_out[527]
  PIN data_out[528]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2164.000 0.000 2164.600 ;
    END
  END data_out[528]
  PIN data_out[529]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2168.000 0.000 2168.600 ;
    END
  END data_out[529]
  PIN data_out[530]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2172.000 0.000 2172.600 ;
    END
  END data_out[530]
  PIN data_out[531]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2176.000 0.000 2176.600 ;
    END
  END data_out[531]
  PIN data_out[532]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2180.000 0.000 2180.600 ;
    END
  END data_out[532]
  PIN data_out[533]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2184.000 0.000 2184.600 ;
    END
  END data_out[533]
  PIN data_out[534]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2188.000 0.000 2188.600 ;
    END
  END data_out[534]
  PIN data_out[535]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2192.000 0.000 2192.600 ;
    END
  END data_out[535]
  PIN data_out[536]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2196.000 0.000 2196.600 ;
    END
  END data_out[536]
  PIN data_out[537]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2200.000 0.000 2200.600 ;
    END
  END data_out[537]
  PIN data_out[538]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2204.000 0.000 2204.600 ;
    END
  END data_out[538]
  PIN data_out[539]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2208.000 0.000 2208.600 ;
    END
  END data_out[539]
  PIN data_out[540]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2212.000 0.000 2212.600 ;
    END
  END data_out[540]
  PIN data_out[541]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2216.000 0.000 2216.600 ;
    END
  END data_out[541]
  PIN data_out[542]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2220.000 0.000 2220.600 ;
    END
  END data_out[542]
  PIN data_out[543]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2224.000 0.000 2224.600 ;
    END
  END data_out[543]
  PIN data_out[544]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2228.000 0.000 2228.600 ;
    END
  END data_out[544]
  PIN data_out[545]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2232.000 0.000 2232.600 ;
    END
  END data_out[545]
  PIN data_out[546]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2236.000 0.000 2236.600 ;
    END
  END data_out[546]
  PIN data_out[547]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2240.000 0.000 2240.600 ;
    END
  END data_out[547]
  PIN data_out[548]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2244.000 0.000 2244.600 ;
    END
  END data_out[548]
  PIN data_out[549]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2248.000 0.000 2248.600 ;
    END
  END data_out[549]
  PIN data_out[550]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2252.000 0.000 2252.600 ;
    END
  END data_out[550]
  PIN data_out[551]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2256.000 0.000 2256.600 ;
    END
  END data_out[551]
  PIN data_out[552]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2260.000 0.000 2260.600 ;
    END
  END data_out[552]
  PIN data_out[553]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2264.000 0.000 2264.600 ;
    END
  END data_out[553]
  PIN data_out[554]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2268.000 0.000 2268.600 ;
    END
  END data_out[554]
  PIN data_out[555]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2272.000 0.000 2272.600 ;
    END
  END data_out[555]
  PIN data_out[556]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2276.000 0.000 2276.600 ;
    END
  END data_out[556]
  PIN data_out[557]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2280.000 0.000 2280.600 ;
    END
  END data_out[557]
  PIN data_out[558]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2284.000 0.000 2284.600 ;
    END
  END data_out[558]
  PIN data_out[559]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2288.000 0.000 2288.600 ;
    END
  END data_out[559]
  PIN data_out[560]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2292.000 0.000 2292.600 ;
    END
  END data_out[560]
  PIN data_out[561]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2296.000 0.000 2296.600 ;
    END
  END data_out[561]
  PIN data_out[562]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2300.000 0.000 2300.600 ;
    END
  END data_out[562]
  PIN data_out[563]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2304.000 0.000 2304.600 ;
    END
  END data_out[563]
  PIN data_out[564]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2308.000 0.000 2308.600 ;
    END
  END data_out[564]
  PIN data_out[565]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2312.000 0.000 2312.600 ;
    END
  END data_out[565]
  PIN data_out[566]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2316.000 0.000 2316.600 ;
    END
  END data_out[566]
  PIN data_out[567]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2320.000 0.000 2320.600 ;
    END
  END data_out[567]
  PIN data_out[568]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2324.000 0.000 2324.600 ;
    END
  END data_out[568]
  PIN data_out[569]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2328.000 0.000 2328.600 ;
    END
  END data_out[569]
  PIN data_out[570]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2332.000 0.000 2332.600 ;
    END
  END data_out[570]
  PIN data_out[571]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2336.000 0.000 2336.600 ;
    END
  END data_out[571]
  PIN data_out[572]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2340.000 0.000 2340.600 ;
    END
  END data_out[572]
  PIN data_out[573]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2344.000 0.000 2344.600 ;
    END
  END data_out[573]
  PIN data_out[574]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2348.000 0.000 2348.600 ;
    END
  END data_out[574]
  PIN data_out[575]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2352.000 0.000 2352.600 ;
    END
  END data_out[575]
  PIN data_out[576]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2356.000 0.000 2356.600 ;
    END
  END data_out[576]
  PIN data_out[577]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2360.000 0.000 2360.600 ;
    END
  END data_out[577]
  PIN data_out[578]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2364.000 0.000 2364.600 ;
    END
  END data_out[578]
  PIN data_out[579]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2368.000 0.000 2368.600 ;
    END
  END data_out[579]
  PIN data_out[580]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2372.000 0.000 2372.600 ;
    END
  END data_out[580]
  PIN data_out[581]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2376.000 0.000 2376.600 ;
    END
  END data_out[581]
  PIN data_out[582]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2380.000 0.000 2380.600 ;
    END
  END data_out[582]
  PIN data_out[583]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2384.000 0.000 2384.600 ;
    END
  END data_out[583]
  PIN data_out[584]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2388.000 0.000 2388.600 ;
    END
  END data_out[584]
  PIN data_out[585]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2392.000 0.000 2392.600 ;
    END
  END data_out[585]
  PIN data_out[586]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2396.000 0.000 2396.600 ;
    END
  END data_out[586]
  PIN data_out[587]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2400.000 0.000 2400.600 ;
    END
  END data_out[587]
  PIN data_out[588]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2404.000 0.000 2404.600 ;
    END
  END data_out[588]
  PIN data_out[589]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2408.000 0.000 2408.600 ;
    END
  END data_out[589]
  PIN data_out[590]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2412.000 0.000 2412.600 ;
    END
  END data_out[590]
  PIN data_out[591]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2416.000 0.000 2416.600 ;
    END
  END data_out[591]
  PIN data_out[592]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2420.000 0.000 2420.600 ;
    END
  END data_out[592]
  PIN data_out[593]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2424.000 0.000 2424.600 ;
    END
  END data_out[593]
  PIN data_out[594]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2428.000 0.000 2428.600 ;
    END
  END data_out[594]
  PIN data_out[595]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2432.000 0.000 2432.600 ;
    END
  END data_out[595]
  PIN data_out[596]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2436.000 0.000 2436.600 ;
    END
  END data_out[596]
  PIN data_out[597]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2440.000 0.000 2440.600 ;
    END
  END data_out[597]
  PIN data_out[598]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2444.000 0.000 2444.600 ;
    END
  END data_out[598]
  PIN data_out[599]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2448.000 0.000 2448.600 ;
    END
  END data_out[599]
  PIN data_out[600]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2452.000 0.000 2452.600 ;
    END
  END data_out[600]
  PIN data_out[601]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2456.000 0.000 2456.600 ;
    END
  END data_out[601]
  PIN data_out[602]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2460.000 0.000 2460.600 ;
    END
  END data_out[602]
  PIN data_out[603]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2464.000 0.000 2464.600 ;
    END
  END data_out[603]
  PIN data_out[604]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2468.000 0.000 2468.600 ;
    END
  END data_out[604]
  PIN data_out[605]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2472.000 0.000 2472.600 ;
    END
  END data_out[605]
  PIN data_out[606]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2476.000 0.000 2476.600 ;
    END
  END data_out[606]
  PIN data_out[607]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2480.000 0.000 2480.600 ;
    END
  END data_out[607]
  PIN data_out[608]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2484.000 0.000 2484.600 ;
    END
  END data_out[608]
  PIN data_out[609]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2488.000 0.000 2488.600 ;
    END
  END data_out[609]
  PIN data_out[610]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2492.000 0.000 2492.600 ;
    END
  END data_out[610]
  PIN data_out[611]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2496.000 0.000 2496.600 ;
    END
  END data_out[611]
  PIN data_out[612]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2500.000 0.000 2500.600 ;
    END
  END data_out[612]
  PIN data_out[613]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2504.000 0.000 2504.600 ;
    END
  END data_out[613]
  PIN data_out[614]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2508.000 0.000 2508.600 ;
    END
  END data_out[614]
  PIN data_out[615]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2512.000 0.000 2512.600 ;
    END
  END data_out[615]
  PIN data_out[616]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2516.000 0.000 2516.600 ;
    END
  END data_out[616]
  PIN data_out[617]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2520.000 0.000 2520.600 ;
    END
  END data_out[617]
  PIN data_out[618]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2524.000 0.000 2524.600 ;
    END
  END data_out[618]
  PIN data_out[619]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2528.000 0.000 2528.600 ;
    END
  END data_out[619]
  PIN data_out[620]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2532.000 0.000 2532.600 ;
    END
  END data_out[620]
  PIN data_out[621]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2536.000 0.000 2536.600 ;
    END
  END data_out[621]
  PIN data_out[622]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2540.000 0.000 2540.600 ;
    END
  END data_out[622]
  PIN data_out[623]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2544.000 0.000 2544.600 ;
    END
  END data_out[623]
  PIN data_out[624]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2548.000 0.000 2548.600 ;
    END
  END data_out[624]
  PIN data_out[625]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2552.000 0.000 2552.600 ;
    END
  END data_out[625]
  PIN data_out[626]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2556.000 0.000 2556.600 ;
    END
  END data_out[626]
  PIN data_out[627]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2560.000 0.000 2560.600 ;
    END
  END data_out[627]
  PIN data_out[628]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2564.000 0.000 2564.600 ;
    END
  END data_out[628]
  PIN data_out[629]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2568.000 0.000 2568.600 ;
    END
  END data_out[629]
  PIN data_out[630]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2572.000 0.000 2572.600 ;
    END
  END data_out[630]
  PIN data_out[631]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2576.000 0.000 2576.600 ;
    END
  END data_out[631]
  PIN data_out[632]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2580.000 0.000 2580.600 ;
    END
  END data_out[632]
  PIN data_out[633]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2584.000 0.000 2584.600 ;
    END
  END data_out[633]
  PIN data_out[634]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2588.000 0.000 2588.600 ;
    END
  END data_out[634]
  PIN data_out[635]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2592.000 0.000 2592.600 ;
    END
  END data_out[635]
  PIN data_out[636]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2596.000 0.000 2596.600 ;
    END
  END data_out[636]
  PIN data_out[637]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2600.000 0.000 2600.600 ;
    END
  END data_out[637]
  PIN data_out[638]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2604.000 0.000 2604.600 ;
    END
  END data_out[638]
  PIN data_out[639]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2608.000 0.000 2608.600 ;
    END
  END data_out[639]
  PIN data_out[640]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2612.000 0.000 2612.600 ;
    END
  END data_out[640]
  PIN data_out[641]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2616.000 0.000 2616.600 ;
    END
  END data_out[641]
  PIN data_out[642]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2620.000 0.000 2620.600 ;
    END
  END data_out[642]
  PIN data_out[643]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2624.000 0.000 2624.600 ;
    END
  END data_out[643]
  PIN data_out[644]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2628.000 0.000 2628.600 ;
    END
  END data_out[644]
  PIN data_out[645]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2632.000 0.000 2632.600 ;
    END
  END data_out[645]
  PIN data_out[646]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2636.000 0.000 2636.600 ;
    END
  END data_out[646]
  PIN data_out[647]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 2640.000 0.000 2640.600 ;
    END
  END data_out[647]
END tri_512x162_4w_0
END LIBRARY


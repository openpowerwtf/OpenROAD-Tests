VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO toysram_bare_32x32_2r1w
  CLASS BLOCK ;
  FOREIGN toysram_bare_32x32_2r1w ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 150.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.000 0.000 4.600 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 6.000 0.000 6.600 ;
    END
  END GND
  PIN rd0_c_na0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 4.000 104.000 4.600 ;
    END
  END rd0_c_na0
  PIN rd0_c_a0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 6.000 104.000 6.600 ;
    END
  END rd0_c_a0
  PIN rd0_na1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 8.000 104.000 8.600 ;
    END
  END rd0_na1_na2
  PIN rd0_na1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 10.000 104.000 10.600 ;
    END
  END rd0_na1_a2
  PIN rd0_a1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 12.000 104.000 12.600 ;
    END
  END rd0_a1_na2
  PIN rd0_a1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 14.000 104.000 14.600 ;
    END
  END rd0_a1_a2
  PIN rd0_na3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 16.000 104.000 16.600 ;
    END
  END rd0_na3
  PIN rd0_a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 18.000 104.000 18.600 ;
    END
  END rd0_a3
  PIN rd0_na4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 20.000 104.000 20.600 ;
    END
  END rd0_na4
  PIN rd0_a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 22.000 104.000 22.600 ;
    END
  END rd0_a4
  PIN rd1_c_na0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 24.000 104.000 24.600 ;
    END
  END rd1_c_na0
  PIN rd1_c_a0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 26.000 104.000 26.600 ;
    END
  END rd1_c_a0
  PIN rd1_na1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 28.000 104.000 28.600 ;
    END
  END rd1_na1_na2
  PIN rd1_na1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 30.000 104.000 30.600 ;
    END
  END rd1_na1_a2
  PIN rd1_a1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 32.000 104.000 32.600 ;
    END
  END rd1_a1_na2
  PIN rd1_a1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 34.000 104.000 34.600 ;
    END
  END rd1_a1_a2
  PIN rd1_na3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 36.000 104.000 36.600 ;
    END
  END rd1_na3
  PIN rd1_a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 38.000 104.000 38.600 ;
    END
  END rd1_a3
  PIN rd1_na4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 40.000 104.000 40.600 ;
    END
  END rd1_na4
  PIN rd1_a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 42.000 104.000 42.600 ;
    END
  END rd1_a4
  PIN wr0_c_na0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 44.000 104.000 44.600 ;
    END
  END wr0_c_na0
  PIN wr0_c_a0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 46.000 104.000 46.600 ;
    END
  END wr0_c_a0
  PIN wr0_na1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 48.000 104.000 48.600 ;
    END
  END wr0_na1_na2
  PIN wr0_na1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 50.000 104.000 50.600 ;
    END
  END wr0_na1_a2
  PIN wr0_a1_na2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 52.000 104.000 52.600 ;
    END
  END wr0_a1_na2
  PIN wr0_a1_a2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 54.000 104.000 54.600 ;
    END
  END wr0_a1_a2
  PIN wr0_na3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 56.000 104.000 56.600 ;
    END
  END wr0_na3
  PIN wr0_a3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 58.000 104.000 58.600 ;
    END
  END wr0_a3
  PIN wr0_na4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 60.000 104.000 60.600 ;
    END
  END wr0_na4
  PIN wr0_a4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 62.000 104.000 62.600 ;
    END
  END wr0_a4
  PIN rd0_dat[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.000 0.000 8.600 ;
    END
  END rd0_dat[31]
  PIN rd0_dat[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 10.000 0.000 10.600 ;
    END
  END rd0_dat[30]
  PIN rd0_dat[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.000 0.000 12.600 ;
    END
  END rd0_dat[29]
  PIN rd0_dat[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 14.000 0.000 14.600 ;
    END
  END rd0_dat[28]
  PIN rd0_dat[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 16.000 0.000 16.600 ;
    END
  END rd0_dat[27]
  PIN rd0_dat[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 18.000 0.000 18.600 ;
    END
  END rd0_dat[26]
  PIN rd0_dat[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 20.000 0.000 20.600 ;
    END
  END rd0_dat[25]
  PIN rd0_dat[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 22.000 0.000 22.600 ;
    END
  END rd0_dat[24]
  PIN rd0_dat[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 24.000 0.000 24.600 ;
    END
  END rd0_dat[23]
  PIN rd0_dat[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 26.000 0.000 26.600 ;
    END
  END rd0_dat[22]
  PIN rd0_dat[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 28.000 0.000 28.600 ;
    END
  END rd0_dat[21]
  PIN rd0_dat[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 30.000 0.000 30.600 ;
    END
  END rd0_dat[20]
  PIN rd0_dat[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 0.000 32.600 ;
    END
  END rd0_dat[19]
  PIN rd0_dat[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 34.000 0.000 34.600 ;
    END
  END rd0_dat[18]
  PIN rd0_dat[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.000 0.000 36.600 ;
    END
  END rd0_dat[17]
  PIN rd0_dat[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 38.000 0.000 38.600 ;
    END
  END rd0_dat[16]
  PIN rd0_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.000 0.000 40.600 ;
    END
  END rd0_dat[15]
  PIN rd0_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 42.000 0.000 42.600 ;
    END
  END rd0_dat[14]
  PIN rd0_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.000 0.000 44.600 ;
    END
  END rd0_dat[13]
  PIN rd0_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 46.000 0.000 46.600 ;
    END
  END rd0_dat[12]
  PIN rd0_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.000 0.000 48.600 ;
    END
  END rd0_dat[11]
  PIN rd0_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 50.000 0.000 50.600 ;
    END
  END rd0_dat[10]
  PIN rd0_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 52.000 0.000 52.600 ;
    END
  END rd0_dat[9]
  PIN rd0_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 54.000 0.000 54.600 ;
    END
  END rd0_dat[8]
  PIN rd0_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 56.000 0.000 56.600 ;
    END
  END rd0_dat[7]
  PIN rd0_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 58.000 0.000 58.600 ;
    END
  END rd0_dat[6]
  PIN rd0_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 60.000 0.000 60.600 ;
    END
  END rd0_dat[5]
  PIN rd0_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 62.000 0.000 62.600 ;
    END
  END rd0_dat[4]
  PIN rd0_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 64.000 0.000 64.600 ;
    END
  END rd0_dat[3]
  PIN rd0_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 66.000 0.000 66.600 ;
    END
  END rd0_dat[2]
  PIN rd0_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.000 0.000 68.600 ;
    END
  END rd0_dat[1]
  PIN rd0_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 70.000 0.000 70.600 ;
    END
  END rd0_dat[0]
  PIN rd1_dat[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.000 0.000 72.600 ;
    END
  END rd1_dat[31]
  PIN rd1_dat[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 74.000 0.000 74.600 ;
    END
  END rd1_dat[30]
  PIN rd1_dat[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.000 0.000 76.600 ;
    END
  END rd1_dat[29]
  PIN rd1_dat[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 78.000 0.000 78.600 ;
    END
  END rd1_dat[28]
  PIN rd1_dat[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.000 0.000 80.600 ;
    END
  END rd1_dat[27]
  PIN rd1_dat[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 82.000 0.000 82.600 ;
    END
  END rd1_dat[26]
  PIN rd1_dat[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.000 0.000 84.600 ;
    END
  END rd1_dat[25]
  PIN rd1_dat[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 86.000 0.000 86.600 ;
    END
  END rd1_dat[24]
  PIN rd1_dat[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.000 0.000 88.600 ;
    END
  END rd1_dat[23]
  PIN rd1_dat[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 90.000 0.000 90.600 ;
    END
  END rd1_dat[22]
  PIN rd1_dat[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.000 0.000 92.600 ;
    END
  END rd1_dat[21]
  PIN rd1_dat[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 94.000 0.000 94.600 ;
    END
  END rd1_dat[20]
  PIN rd1_dat[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.000 0.000 96.600 ;
    END
  END rd1_dat[19]
  PIN rd1_dat[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 98.000 0.000 98.600 ;
    END
  END rd1_dat[18]
  PIN rd1_dat[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.000 0.000 100.600 ;
    END
  END rd1_dat[17]
  PIN rd1_dat[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 102.000 0.000 102.600 ;
    END
  END rd1_dat[16]
  PIN rd1_dat[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.000 0.000 104.600 ;
    END
  END rd1_dat[15]
  PIN rd1_dat[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 106.000 0.000 106.600 ;
    END
  END rd1_dat[14]
  PIN rd1_dat[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.000 0.000 108.600 ;
    END
  END rd1_dat[13]
  PIN rd1_dat[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 110.000 0.000 110.600 ;
    END
  END rd1_dat[12]
  PIN rd1_dat[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.000 0.000 112.600 ;
    END
  END rd1_dat[11]
  PIN rd1_dat[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 114.000 0.000 114.600 ;
    END
  END rd1_dat[10]
  PIN rd1_dat[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 116.000 0.000 116.600 ;
    END
  END rd1_dat[9]
  PIN rd1_dat[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 118.000 0.000 118.600 ;
    END
  END rd1_dat[8]
  PIN rd1_dat[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 120.000 0.000 120.600 ;
    END
  END rd1_dat[7]
  PIN rd1_dat[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 122.000 0.000 122.600 ;
    END
  END rd1_dat[6]
  PIN rd1_dat[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 124.000 0.000 124.600 ;
    END
  END rd1_dat[5]
  PIN rd1_dat[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 126.000 0.000 126.600 ;
    END
  END rd1_dat[4]
  PIN rd1_dat[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 128.000 0.000 128.600 ;
    END
  END rd1_dat[3]
  PIN rd1_dat[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 130.000 0.000 130.600 ;
    END
  END rd1_dat[2]
  PIN rd1_dat[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 132.000 0.000 132.600 ;
    END
  END rd1_dat[1]
  PIN rd1_dat[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 134.000 0.000 134.600 ;
    END
  END rd1_dat[0]
  PIN wr0_dat[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 64.000 104.000 64.600 ;
    END
  END wr0_dat[31]
  PIN wr0_dat[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 66.000 104.000 66.600 ;
    END
  END wr0_dat[30]
  PIN wr0_dat[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 68.000 104.000 68.600 ;
    END
  END wr0_dat[29]
  PIN wr0_dat[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 70.000 104.000 70.600 ;
    END
  END wr0_dat[28]
  PIN wr0_dat[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 72.000 104.000 72.600 ;
    END
  END wr0_dat[27]
  PIN wr0_dat[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 74.000 104.000 74.600 ;
    END
  END wr0_dat[26]
  PIN wr0_dat[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 76.000 104.000 76.600 ;
    END
  END wr0_dat[25]
  PIN wr0_dat[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 78.000 104.000 78.600 ;
    END
  END wr0_dat[24]
  PIN wr0_dat[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 80.000 104.000 80.600 ;
    END
  END wr0_dat[23]
  PIN wr0_dat[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 82.000 104.000 82.600 ;
    END
  END wr0_dat[22]
  PIN wr0_dat[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 84.000 104.000 84.600 ;
    END
  END wr0_dat[21]
  PIN wr0_dat[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 86.000 104.000 86.600 ;
    END
  END wr0_dat[20]
  PIN wr0_dat[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 88.000 104.000 88.600 ;
    END
  END wr0_dat[19]
  PIN wr0_dat[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 90.000 104.000 90.600 ;
    END
  END wr0_dat[18]
  PIN wr0_dat[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 92.000 104.000 92.600 ;
    END
  END wr0_dat[17]
  PIN wr0_dat[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 94.000 104.000 94.600 ;
    END
  END wr0_dat[16]
  PIN wr0_dat[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 96.000 104.000 96.600 ;
    END
  END wr0_dat[15]
  PIN wr0_dat[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 98.000 104.000 98.600 ;
    END
  END wr0_dat[14]
  PIN wr0_dat[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 100.000 104.000 100.600 ;
    END
  END wr0_dat[13]
  PIN wr0_dat[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 102.000 104.000 102.600 ;
    END
  END wr0_dat[12]
  PIN wr0_dat[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 104.000 104.000 104.600 ;
    END
  END wr0_dat[11]
  PIN wr0_dat[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 106.000 104.000 106.600 ;
    END
  END wr0_dat[10]
  PIN wr0_dat[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 108.000 104.000 108.600 ;
    END
  END wr0_dat[9]
  PIN wr0_dat[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 110.000 104.000 110.600 ;
    END
  END wr0_dat[8]
  PIN wr0_dat[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 112.000 104.000 112.600 ;
    END
  END wr0_dat[7]
  PIN wr0_dat[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 114.000 104.000 114.600 ;
    END
  END wr0_dat[6]
  PIN wr0_dat[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 116.000 104.000 116.600 ;
    END
  END wr0_dat[5]
  PIN wr0_dat[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 118.000 104.000 118.600 ;
    END
  END wr0_dat[4]
  PIN wr0_dat[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 120.000 104.000 120.600 ;
    END
  END wr0_dat[3]
  PIN wr0_dat[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 122.000 104.000 122.600 ;
    END
  END wr0_dat[2]
  PIN wr0_dat[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 124.000 104.000 124.600 ;
    END
  END wr0_dat[1]
  PIN wr0_dat[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.000 126.000 104.000 126.600 ;
    END
  END wr0_dat[0]
END toysram_bare_32x32_2r1w
END LIBRARY


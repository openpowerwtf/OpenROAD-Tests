VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tri_fu_mul
  CLASS BLOCK ;
  FOREIGN tri_fu_mul ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 900.000 ;
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 4.000 0.000 4.600 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 8.000 0.000 8.600 ;
    END
  END gnd
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 4.000 254.000 4.600 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 8.000 254.000 8.600 ;
    END
  END rst
  PIN clkoff_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 12.000 254.000 12.600 ;
    END
  END clkoff_b
  PIN act_dis
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 16.000 254.000 16.600 ;
    END
  END act_dis
  PIN flush
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 20.000 254.000 20.600 ;
    END
  END flush
  PIN delay_lclkr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 24.000 254.000 24.600 ;
    END
  END delay_lclkr
  PIN mpw1_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 28.000 254.000 28.600 ;
    END
  END mpw1_b
  PIN mpw2_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 32.000 254.000 32.600 ;
    END
  END mpw2_b
  PIN sg_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 36.000 254.000 36.600 ;
    END
  END sg_1
  PIN thold_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 40.000 254.000 40.600 ;
    END
  END thold_1
  PIN fpu_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 44.000 254.000 44.600 ;
    END
  END fpu_enable
  PIN f_mul_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 48.000 254.000 48.600 ;
    END
  END f_mul_si
  PIN f_mul_so
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 12.000 0.000 12.600 ;
    END
  END f_mul_so
  PIN ex2_act
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 52.000 254.000 52.600 ;
    END
  END ex2_act
  PIN f_fmt_ex2_a_frac[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 56.000 254.000 56.600 ;
    END
  END f_fmt_ex2_a_frac[0]
  PIN f_fmt_ex2_a_frac[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 60.000 254.000 60.600 ;
    END
  END f_fmt_ex2_a_frac[1]
  PIN f_fmt_ex2_a_frac[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 64.000 254.000 64.600 ;
    END
  END f_fmt_ex2_a_frac[2]
  PIN f_fmt_ex2_a_frac[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 68.000 254.000 68.600 ;
    END
  END f_fmt_ex2_a_frac[3]
  PIN f_fmt_ex2_a_frac[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 72.000 254.000 72.600 ;
    END
  END f_fmt_ex2_a_frac[4]
  PIN f_fmt_ex2_a_frac[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 76.000 254.000 76.600 ;
    END
  END f_fmt_ex2_a_frac[5]
  PIN f_fmt_ex2_a_frac[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 80.000 254.000 80.600 ;
    END
  END f_fmt_ex2_a_frac[6]
  PIN f_fmt_ex2_a_frac[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 84.000 254.000 84.600 ;
    END
  END f_fmt_ex2_a_frac[7]
  PIN f_fmt_ex2_a_frac[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 88.000 254.000 88.600 ;
    END
  END f_fmt_ex2_a_frac[8]
  PIN f_fmt_ex2_a_frac[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 92.000 254.000 92.600 ;
    END
  END f_fmt_ex2_a_frac[9]
  PIN f_fmt_ex2_a_frac[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 96.000 254.000 96.600 ;
    END
  END f_fmt_ex2_a_frac[10]
  PIN f_fmt_ex2_a_frac[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 100.000 254.000 100.600 ;
    END
  END f_fmt_ex2_a_frac[11]
  PIN f_fmt_ex2_a_frac[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 104.000 254.000 104.600 ;
    END
  END f_fmt_ex2_a_frac[12]
  PIN f_fmt_ex2_a_frac[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 108.000 254.000 108.600 ;
    END
  END f_fmt_ex2_a_frac[13]
  PIN f_fmt_ex2_a_frac[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 112.000 254.000 112.600 ;
    END
  END f_fmt_ex2_a_frac[14]
  PIN f_fmt_ex2_a_frac[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 116.000 254.000 116.600 ;
    END
  END f_fmt_ex2_a_frac[15]
  PIN f_fmt_ex2_a_frac[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 120.000 254.000 120.600 ;
    END
  END f_fmt_ex2_a_frac[16]
  PIN f_fmt_ex2_a_frac[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 124.000 254.000 124.600 ;
    END
  END f_fmt_ex2_a_frac[17]
  PIN f_fmt_ex2_a_frac[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 128.000 254.000 128.600 ;
    END
  END f_fmt_ex2_a_frac[18]
  PIN f_fmt_ex2_a_frac[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 132.000 254.000 132.600 ;
    END
  END f_fmt_ex2_a_frac[19]
  PIN f_fmt_ex2_a_frac[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 136.000 254.000 136.600 ;
    END
  END f_fmt_ex2_a_frac[20]
  PIN f_fmt_ex2_a_frac[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 140.000 254.000 140.600 ;
    END
  END f_fmt_ex2_a_frac[21]
  PIN f_fmt_ex2_a_frac[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 144.000 254.000 144.600 ;
    END
  END f_fmt_ex2_a_frac[22]
  PIN f_fmt_ex2_a_frac[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 148.000 254.000 148.600 ;
    END
  END f_fmt_ex2_a_frac[23]
  PIN f_fmt_ex2_a_frac[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 152.000 254.000 152.600 ;
    END
  END f_fmt_ex2_a_frac[24]
  PIN f_fmt_ex2_a_frac[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 156.000 254.000 156.600 ;
    END
  END f_fmt_ex2_a_frac[25]
  PIN f_fmt_ex2_a_frac[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 160.000 254.000 160.600 ;
    END
  END f_fmt_ex2_a_frac[26]
  PIN f_fmt_ex2_a_frac[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 164.000 254.000 164.600 ;
    END
  END f_fmt_ex2_a_frac[27]
  PIN f_fmt_ex2_a_frac[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 168.000 254.000 168.600 ;
    END
  END f_fmt_ex2_a_frac[28]
  PIN f_fmt_ex2_a_frac[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 172.000 254.000 172.600 ;
    END
  END f_fmt_ex2_a_frac[29]
  PIN f_fmt_ex2_a_frac[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 176.000 254.000 176.600 ;
    END
  END f_fmt_ex2_a_frac[30]
  PIN f_fmt_ex2_a_frac[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 180.000 254.000 180.600 ;
    END
  END f_fmt_ex2_a_frac[31]
  PIN f_fmt_ex2_a_frac[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 184.000 254.000 184.600 ;
    END
  END f_fmt_ex2_a_frac[32]
  PIN f_fmt_ex2_a_frac[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 188.000 254.000 188.600 ;
    END
  END f_fmt_ex2_a_frac[33]
  PIN f_fmt_ex2_a_frac[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 192.000 254.000 192.600 ;
    END
  END f_fmt_ex2_a_frac[34]
  PIN f_fmt_ex2_a_frac[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 196.000 254.000 196.600 ;
    END
  END f_fmt_ex2_a_frac[35]
  PIN f_fmt_ex2_a_frac[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 200.000 254.000 200.600 ;
    END
  END f_fmt_ex2_a_frac[36]
  PIN f_fmt_ex2_a_frac[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 204.000 254.000 204.600 ;
    END
  END f_fmt_ex2_a_frac[37]
  PIN f_fmt_ex2_a_frac[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 208.000 254.000 208.600 ;
    END
  END f_fmt_ex2_a_frac[38]
  PIN f_fmt_ex2_a_frac[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 212.000 254.000 212.600 ;
    END
  END f_fmt_ex2_a_frac[39]
  PIN f_fmt_ex2_a_frac[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 216.000 254.000 216.600 ;
    END
  END f_fmt_ex2_a_frac[40]
  PIN f_fmt_ex2_a_frac[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 220.000 254.000 220.600 ;
    END
  END f_fmt_ex2_a_frac[41]
  PIN f_fmt_ex2_a_frac[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 224.000 254.000 224.600 ;
    END
  END f_fmt_ex2_a_frac[42]
  PIN f_fmt_ex2_a_frac[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 228.000 254.000 228.600 ;
    END
  END f_fmt_ex2_a_frac[43]
  PIN f_fmt_ex2_a_frac[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 232.000 254.000 232.600 ;
    END
  END f_fmt_ex2_a_frac[44]
  PIN f_fmt_ex2_a_frac[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 236.000 254.000 236.600 ;
    END
  END f_fmt_ex2_a_frac[45]
  PIN f_fmt_ex2_a_frac[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 240.000 254.000 240.600 ;
    END
  END f_fmt_ex2_a_frac[46]
  PIN f_fmt_ex2_a_frac[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 244.000 254.000 244.600 ;
    END
  END f_fmt_ex2_a_frac[47]
  PIN f_fmt_ex2_a_frac[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 248.000 254.000 248.600 ;
    END
  END f_fmt_ex2_a_frac[48]
  PIN f_fmt_ex2_a_frac[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 252.000 254.000 252.600 ;
    END
  END f_fmt_ex2_a_frac[49]
  PIN f_fmt_ex2_a_frac[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 256.000 254.000 256.600 ;
    END
  END f_fmt_ex2_a_frac[50]
  PIN f_fmt_ex2_a_frac[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 260.000 254.000 260.600 ;
    END
  END f_fmt_ex2_a_frac[51]
  PIN f_fmt_ex2_a_frac[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 264.000 254.000 264.600 ;
    END
  END f_fmt_ex2_a_frac[52]
  PIN f_fmt_ex2_a_frac_17
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 268.000 254.000 268.600 ;
    END
  END f_fmt_ex2_a_frac_17
  PIN f_fmt_ex2_a_frac_35
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 272.000 254.000 272.600 ;
    END
  END f_fmt_ex2_a_frac_35
  PIN f_fmt_ex2_c_frac[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 276.000 254.000 276.600 ;
    END
  END f_fmt_ex2_c_frac[0]
  PIN f_fmt_ex2_c_frac[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 280.000 254.000 280.600 ;
    END
  END f_fmt_ex2_c_frac[1]
  PIN f_fmt_ex2_c_frac[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 284.000 254.000 284.600 ;
    END
  END f_fmt_ex2_c_frac[2]
  PIN f_fmt_ex2_c_frac[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 288.000 254.000 288.600 ;
    END
  END f_fmt_ex2_c_frac[3]
  PIN f_fmt_ex2_c_frac[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 292.000 254.000 292.600 ;
    END
  END f_fmt_ex2_c_frac[4]
  PIN f_fmt_ex2_c_frac[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 296.000 254.000 296.600 ;
    END
  END f_fmt_ex2_c_frac[5]
  PIN f_fmt_ex2_c_frac[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 300.000 254.000 300.600 ;
    END
  END f_fmt_ex2_c_frac[6]
  PIN f_fmt_ex2_c_frac[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 304.000 254.000 304.600 ;
    END
  END f_fmt_ex2_c_frac[7]
  PIN f_fmt_ex2_c_frac[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 308.000 254.000 308.600 ;
    END
  END f_fmt_ex2_c_frac[8]
  PIN f_fmt_ex2_c_frac[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 312.000 254.000 312.600 ;
    END
  END f_fmt_ex2_c_frac[9]
  PIN f_fmt_ex2_c_frac[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 316.000 254.000 316.600 ;
    END
  END f_fmt_ex2_c_frac[10]
  PIN f_fmt_ex2_c_frac[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 320.000 254.000 320.600 ;
    END
  END f_fmt_ex2_c_frac[11]
  PIN f_fmt_ex2_c_frac[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 324.000 254.000 324.600 ;
    END
  END f_fmt_ex2_c_frac[12]
  PIN f_fmt_ex2_c_frac[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 328.000 254.000 328.600 ;
    END
  END f_fmt_ex2_c_frac[13]
  PIN f_fmt_ex2_c_frac[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 332.000 254.000 332.600 ;
    END
  END f_fmt_ex2_c_frac[14]
  PIN f_fmt_ex2_c_frac[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 336.000 254.000 336.600 ;
    END
  END f_fmt_ex2_c_frac[15]
  PIN f_fmt_ex2_c_frac[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 340.000 254.000 340.600 ;
    END
  END f_fmt_ex2_c_frac[16]
  PIN f_fmt_ex2_c_frac[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 344.000 254.000 344.600 ;
    END
  END f_fmt_ex2_c_frac[17]
  PIN f_fmt_ex2_c_frac[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 348.000 254.000 348.600 ;
    END
  END f_fmt_ex2_c_frac[18]
  PIN f_fmt_ex2_c_frac[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 352.000 254.000 352.600 ;
    END
  END f_fmt_ex2_c_frac[19]
  PIN f_fmt_ex2_c_frac[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 356.000 254.000 356.600 ;
    END
  END f_fmt_ex2_c_frac[20]
  PIN f_fmt_ex2_c_frac[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 360.000 254.000 360.600 ;
    END
  END f_fmt_ex2_c_frac[21]
  PIN f_fmt_ex2_c_frac[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 364.000 254.000 364.600 ;
    END
  END f_fmt_ex2_c_frac[22]
  PIN f_fmt_ex2_c_frac[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 368.000 254.000 368.600 ;
    END
  END f_fmt_ex2_c_frac[23]
  PIN f_fmt_ex2_c_frac[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 372.000 254.000 372.600 ;
    END
  END f_fmt_ex2_c_frac[24]
  PIN f_fmt_ex2_c_frac[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 376.000 254.000 376.600 ;
    END
  END f_fmt_ex2_c_frac[25]
  PIN f_fmt_ex2_c_frac[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 380.000 254.000 380.600 ;
    END
  END f_fmt_ex2_c_frac[26]
  PIN f_fmt_ex2_c_frac[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 384.000 254.000 384.600 ;
    END
  END f_fmt_ex2_c_frac[27]
  PIN f_fmt_ex2_c_frac[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 388.000 254.000 388.600 ;
    END
  END f_fmt_ex2_c_frac[28]
  PIN f_fmt_ex2_c_frac[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 392.000 254.000 392.600 ;
    END
  END f_fmt_ex2_c_frac[29]
  PIN f_fmt_ex2_c_frac[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 396.000 254.000 396.600 ;
    END
  END f_fmt_ex2_c_frac[30]
  PIN f_fmt_ex2_c_frac[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 400.000 254.000 400.600 ;
    END
  END f_fmt_ex2_c_frac[31]
  PIN f_fmt_ex2_c_frac[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 404.000 254.000 404.600 ;
    END
  END f_fmt_ex2_c_frac[32]
  PIN f_fmt_ex2_c_frac[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 408.000 254.000 408.600 ;
    END
  END f_fmt_ex2_c_frac[33]
  PIN f_fmt_ex2_c_frac[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 412.000 254.000 412.600 ;
    END
  END f_fmt_ex2_c_frac[34]
  PIN f_fmt_ex2_c_frac[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 416.000 254.000 416.600 ;
    END
  END f_fmt_ex2_c_frac[35]
  PIN f_fmt_ex2_c_frac[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 420.000 254.000 420.600 ;
    END
  END f_fmt_ex2_c_frac[36]
  PIN f_fmt_ex2_c_frac[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 424.000 254.000 424.600 ;
    END
  END f_fmt_ex2_c_frac[37]
  PIN f_fmt_ex2_c_frac[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 428.000 254.000 428.600 ;
    END
  END f_fmt_ex2_c_frac[38]
  PIN f_fmt_ex2_c_frac[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 432.000 254.000 432.600 ;
    END
  END f_fmt_ex2_c_frac[39]
  PIN f_fmt_ex2_c_frac[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 436.000 254.000 436.600 ;
    END
  END f_fmt_ex2_c_frac[40]
  PIN f_fmt_ex2_c_frac[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 440.000 254.000 440.600 ;
    END
  END f_fmt_ex2_c_frac[41]
  PIN f_fmt_ex2_c_frac[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 444.000 254.000 444.600 ;
    END
  END f_fmt_ex2_c_frac[42]
  PIN f_fmt_ex2_c_frac[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 448.000 254.000 448.600 ;
    END
  END f_fmt_ex2_c_frac[43]
  PIN f_fmt_ex2_c_frac[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 452.000 254.000 452.600 ;
    END
  END f_fmt_ex2_c_frac[44]
  PIN f_fmt_ex2_c_frac[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 456.000 254.000 456.600 ;
    END
  END f_fmt_ex2_c_frac[45]
  PIN f_fmt_ex2_c_frac[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 460.000 254.000 460.600 ;
    END
  END f_fmt_ex2_c_frac[46]
  PIN f_fmt_ex2_c_frac[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 464.000 254.000 464.600 ;
    END
  END f_fmt_ex2_c_frac[47]
  PIN f_fmt_ex2_c_frac[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 468.000 254.000 468.600 ;
    END
  END f_fmt_ex2_c_frac[48]
  PIN f_fmt_ex2_c_frac[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 472.000 254.000 472.600 ;
    END
  END f_fmt_ex2_c_frac[49]
  PIN f_fmt_ex2_c_frac[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 476.000 254.000 476.600 ;
    END
  END f_fmt_ex2_c_frac[50]
  PIN f_fmt_ex2_c_frac[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 480.000 254.000 480.600 ;
    END
  END f_fmt_ex2_c_frac[51]
  PIN f_fmt_ex2_c_frac[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 484.000 254.000 484.600 ;
    END
  END f_fmt_ex2_c_frac[52]
  PIN f_fmt_ex2_c_frac[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.000 488.000 254.000 488.600 ;
    END
  END f_fmt_ex2_c_frac[53]
  PIN f_mul_ex3_sum[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 16.000 0.000 16.600 ;
    END
  END f_mul_ex3_sum[1]
  PIN f_mul_ex3_sum[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 20.000 0.000 20.600 ;
    END
  END f_mul_ex3_sum[2]
  PIN f_mul_ex3_sum[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 24.000 0.000 24.600 ;
    END
  END f_mul_ex3_sum[3]
  PIN f_mul_ex3_sum[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 28.000 0.000 28.600 ;
    END
  END f_mul_ex3_sum[4]
  PIN f_mul_ex3_sum[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 32.000 0.000 32.600 ;
    END
  END f_mul_ex3_sum[5]
  PIN f_mul_ex3_sum[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 36.000 0.000 36.600 ;
    END
  END f_mul_ex3_sum[6]
  PIN f_mul_ex3_sum[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 40.000 0.000 40.600 ;
    END
  END f_mul_ex3_sum[7]
  PIN f_mul_ex3_sum[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 44.000 0.000 44.600 ;
    END
  END f_mul_ex3_sum[8]
  PIN f_mul_ex3_sum[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 48.000 0.000 48.600 ;
    END
  END f_mul_ex3_sum[9]
  PIN f_mul_ex3_sum[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 52.000 0.000 52.600 ;
    END
  END f_mul_ex3_sum[10]
  PIN f_mul_ex3_sum[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 56.000 0.000 56.600 ;
    END
  END f_mul_ex3_sum[11]
  PIN f_mul_ex3_sum[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 60.000 0.000 60.600 ;
    END
  END f_mul_ex3_sum[12]
  PIN f_mul_ex3_sum[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 64.000 0.000 64.600 ;
    END
  END f_mul_ex3_sum[13]
  PIN f_mul_ex3_sum[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 68.000 0.000 68.600 ;
    END
  END f_mul_ex3_sum[14]
  PIN f_mul_ex3_sum[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 72.000 0.000 72.600 ;
    END
  END f_mul_ex3_sum[15]
  PIN f_mul_ex3_sum[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 76.000 0.000 76.600 ;
    END
  END f_mul_ex3_sum[16]
  PIN f_mul_ex3_sum[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 80.000 0.000 80.600 ;
    END
  END f_mul_ex3_sum[17]
  PIN f_mul_ex3_sum[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 84.000 0.000 84.600 ;
    END
  END f_mul_ex3_sum[18]
  PIN f_mul_ex3_sum[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 88.000 0.000 88.600 ;
    END
  END f_mul_ex3_sum[19]
  PIN f_mul_ex3_sum[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 92.000 0.000 92.600 ;
    END
  END f_mul_ex3_sum[20]
  PIN f_mul_ex3_sum[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 96.000 0.000 96.600 ;
    END
  END f_mul_ex3_sum[21]
  PIN f_mul_ex3_sum[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 100.000 0.000 100.600 ;
    END
  END f_mul_ex3_sum[22]
  PIN f_mul_ex3_sum[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 104.000 0.000 104.600 ;
    END
  END f_mul_ex3_sum[23]
  PIN f_mul_ex3_sum[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 108.000 0.000 108.600 ;
    END
  END f_mul_ex3_sum[24]
  PIN f_mul_ex3_sum[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 112.000 0.000 112.600 ;
    END
  END f_mul_ex3_sum[25]
  PIN f_mul_ex3_sum[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 116.000 0.000 116.600 ;
    END
  END f_mul_ex3_sum[26]
  PIN f_mul_ex3_sum[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 120.000 0.000 120.600 ;
    END
  END f_mul_ex3_sum[27]
  PIN f_mul_ex3_sum[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 124.000 0.000 124.600 ;
    END
  END f_mul_ex3_sum[28]
  PIN f_mul_ex3_sum[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 128.000 0.000 128.600 ;
    END
  END f_mul_ex3_sum[29]
  PIN f_mul_ex3_sum[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 132.000 0.000 132.600 ;
    END
  END f_mul_ex3_sum[30]
  PIN f_mul_ex3_sum[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 136.000 0.000 136.600 ;
    END
  END f_mul_ex3_sum[31]
  PIN f_mul_ex3_sum[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 140.000 0.000 140.600 ;
    END
  END f_mul_ex3_sum[32]
  PIN f_mul_ex3_sum[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 144.000 0.000 144.600 ;
    END
  END f_mul_ex3_sum[33]
  PIN f_mul_ex3_sum[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 148.000 0.000 148.600 ;
    END
  END f_mul_ex3_sum[34]
  PIN f_mul_ex3_sum[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 152.000 0.000 152.600 ;
    END
  END f_mul_ex3_sum[35]
  PIN f_mul_ex3_sum[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 156.000 0.000 156.600 ;
    END
  END f_mul_ex3_sum[36]
  PIN f_mul_ex3_sum[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 160.000 0.000 160.600 ;
    END
  END f_mul_ex3_sum[37]
  PIN f_mul_ex3_sum[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 164.000 0.000 164.600 ;
    END
  END f_mul_ex3_sum[38]
  PIN f_mul_ex3_sum[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 168.000 0.000 168.600 ;
    END
  END f_mul_ex3_sum[39]
  PIN f_mul_ex3_sum[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 172.000 0.000 172.600 ;
    END
  END f_mul_ex3_sum[40]
  PIN f_mul_ex3_sum[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 176.000 0.000 176.600 ;
    END
  END f_mul_ex3_sum[41]
  PIN f_mul_ex3_sum[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 180.000 0.000 180.600 ;
    END
  END f_mul_ex3_sum[42]
  PIN f_mul_ex3_sum[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 184.000 0.000 184.600 ;
    END
  END f_mul_ex3_sum[43]
  PIN f_mul_ex3_sum[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 188.000 0.000 188.600 ;
    END
  END f_mul_ex3_sum[44]
  PIN f_mul_ex3_sum[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 192.000 0.000 192.600 ;
    END
  END f_mul_ex3_sum[45]
  PIN f_mul_ex3_sum[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 196.000 0.000 196.600 ;
    END
  END f_mul_ex3_sum[46]
  PIN f_mul_ex3_sum[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 200.000 0.000 200.600 ;
    END
  END f_mul_ex3_sum[47]
  PIN f_mul_ex3_sum[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 204.000 0.000 204.600 ;
    END
  END f_mul_ex3_sum[48]
  PIN f_mul_ex3_sum[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 208.000 0.000 208.600 ;
    END
  END f_mul_ex3_sum[49]
  PIN f_mul_ex3_sum[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 212.000 0.000 212.600 ;
    END
  END f_mul_ex3_sum[50]
  PIN f_mul_ex3_sum[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 216.000 0.000 216.600 ;
    END
  END f_mul_ex3_sum[51]
  PIN f_mul_ex3_sum[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 220.000 0.000 220.600 ;
    END
  END f_mul_ex3_sum[52]
  PIN f_mul_ex3_sum[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 224.000 0.000 224.600 ;
    END
  END f_mul_ex3_sum[53]
  PIN f_mul_ex3_sum[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 228.000 0.000 228.600 ;
    END
  END f_mul_ex3_sum[54]
  PIN f_mul_ex3_sum[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 232.000 0.000 232.600 ;
    END
  END f_mul_ex3_sum[55]
  PIN f_mul_ex3_sum[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 236.000 0.000 236.600 ;
    END
  END f_mul_ex3_sum[56]
  PIN f_mul_ex3_sum[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 240.000 0.000 240.600 ;
    END
  END f_mul_ex3_sum[57]
  PIN f_mul_ex3_sum[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 244.000 0.000 244.600 ;
    END
  END f_mul_ex3_sum[58]
  PIN f_mul_ex3_sum[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 248.000 0.000 248.600 ;
    END
  END f_mul_ex3_sum[59]
  PIN f_mul_ex3_sum[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 252.000 0.000 252.600 ;
    END
  END f_mul_ex3_sum[60]
  PIN f_mul_ex3_sum[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 256.000 0.000 256.600 ;
    END
  END f_mul_ex3_sum[61]
  PIN f_mul_ex3_sum[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 260.000 0.000 260.600 ;
    END
  END f_mul_ex3_sum[62]
  PIN f_mul_ex3_sum[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 264.000 0.000 264.600 ;
    END
  END f_mul_ex3_sum[63]
  PIN f_mul_ex3_sum[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 268.000 0.000 268.600 ;
    END
  END f_mul_ex3_sum[64]
  PIN f_mul_ex3_sum[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 272.000 0.000 272.600 ;
    END
  END f_mul_ex3_sum[65]
  PIN f_mul_ex3_sum[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 276.000 0.000 276.600 ;
    END
  END f_mul_ex3_sum[66]
  PIN f_mul_ex3_sum[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 280.000 0.000 280.600 ;
    END
  END f_mul_ex3_sum[67]
  PIN f_mul_ex3_sum[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 284.000 0.000 284.600 ;
    END
  END f_mul_ex3_sum[68]
  PIN f_mul_ex3_sum[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 288.000 0.000 288.600 ;
    END
  END f_mul_ex3_sum[69]
  PIN f_mul_ex3_sum[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 292.000 0.000 292.600 ;
    END
  END f_mul_ex3_sum[70]
  PIN f_mul_ex3_sum[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 296.000 0.000 296.600 ;
    END
  END f_mul_ex3_sum[71]
  PIN f_mul_ex3_sum[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 300.000 0.000 300.600 ;
    END
  END f_mul_ex3_sum[72]
  PIN f_mul_ex3_sum[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 304.000 0.000 304.600 ;
    END
  END f_mul_ex3_sum[73]
  PIN f_mul_ex3_sum[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 308.000 0.000 308.600 ;
    END
  END f_mul_ex3_sum[74]
  PIN f_mul_ex3_sum[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 312.000 0.000 312.600 ;
    END
  END f_mul_ex3_sum[75]
  PIN f_mul_ex3_sum[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 316.000 0.000 316.600 ;
    END
  END f_mul_ex3_sum[76]
  PIN f_mul_ex3_sum[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 320.000 0.000 320.600 ;
    END
  END f_mul_ex3_sum[77]
  PIN f_mul_ex3_sum[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 324.000 0.000 324.600 ;
    END
  END f_mul_ex3_sum[78]
  PIN f_mul_ex3_sum[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 328.000 0.000 328.600 ;
    END
  END f_mul_ex3_sum[79]
  PIN f_mul_ex3_sum[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 332.000 0.000 332.600 ;
    END
  END f_mul_ex3_sum[80]
  PIN f_mul_ex3_sum[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 336.000 0.000 336.600 ;
    END
  END f_mul_ex3_sum[81]
  PIN f_mul_ex3_sum[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 340.000 0.000 340.600 ;
    END
  END f_mul_ex3_sum[82]
  PIN f_mul_ex3_sum[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 344.000 0.000 344.600 ;
    END
  END f_mul_ex3_sum[83]
  PIN f_mul_ex3_sum[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 348.000 0.000 348.600 ;
    END
  END f_mul_ex3_sum[84]
  PIN f_mul_ex3_sum[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 352.000 0.000 352.600 ;
    END
  END f_mul_ex3_sum[85]
  PIN f_mul_ex3_sum[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 356.000 0.000 356.600 ;
    END
  END f_mul_ex3_sum[86]
  PIN f_mul_ex3_sum[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 360.000 0.000 360.600 ;
    END
  END f_mul_ex3_sum[87]
  PIN f_mul_ex3_sum[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 364.000 0.000 364.600 ;
    END
  END f_mul_ex3_sum[88]
  PIN f_mul_ex3_sum[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 368.000 0.000 368.600 ;
    END
  END f_mul_ex3_sum[89]
  PIN f_mul_ex3_sum[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 372.000 0.000 372.600 ;
    END
  END f_mul_ex3_sum[90]
  PIN f_mul_ex3_sum[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 376.000 0.000 376.600 ;
    END
  END f_mul_ex3_sum[91]
  PIN f_mul_ex3_sum[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 380.000 0.000 380.600 ;
    END
  END f_mul_ex3_sum[92]
  PIN f_mul_ex3_sum[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 384.000 0.000 384.600 ;
    END
  END f_mul_ex3_sum[93]
  PIN f_mul_ex3_sum[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 388.000 0.000 388.600 ;
    END
  END f_mul_ex3_sum[94]
  PIN f_mul_ex3_sum[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 392.000 0.000 392.600 ;
    END
  END f_mul_ex3_sum[95]
  PIN f_mul_ex3_sum[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 396.000 0.000 396.600 ;
    END
  END f_mul_ex3_sum[96]
  PIN f_mul_ex3_sum[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 400.000 0.000 400.600 ;
    END
  END f_mul_ex3_sum[97]
  PIN f_mul_ex3_sum[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 404.000 0.000 404.600 ;
    END
  END f_mul_ex3_sum[98]
  PIN f_mul_ex3_sum[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 408.000 0.000 408.600 ;
    END
  END f_mul_ex3_sum[99]
  PIN f_mul_ex3_sum[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 412.000 0.000 412.600 ;
    END
  END f_mul_ex3_sum[100]
  PIN f_mul_ex3_sum[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 416.000 0.000 416.600 ;
    END
  END f_mul_ex3_sum[101]
  PIN f_mul_ex3_sum[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 420.000 0.000 420.600 ;
    END
  END f_mul_ex3_sum[102]
  PIN f_mul_ex3_sum[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 424.000 0.000 424.600 ;
    END
  END f_mul_ex3_sum[103]
  PIN f_mul_ex3_sum[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 428.000 0.000 428.600 ;
    END
  END f_mul_ex3_sum[104]
  PIN f_mul_ex3_sum[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 432.000 0.000 432.600 ;
    END
  END f_mul_ex3_sum[105]
  PIN f_mul_ex3_sum[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 436.000 0.000 436.600 ;
    END
  END f_mul_ex3_sum[106]
  PIN f_mul_ex3_sum[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 440.000 0.000 440.600 ;
    END
  END f_mul_ex3_sum[107]
  PIN f_mul_ex3_sum[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 444.000 0.000 444.600 ;
    END
  END f_mul_ex3_sum[108]
  PIN f_mul_ex3_car[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 448.000 0.000 448.600 ;
    END
  END f_mul_ex3_car[1]
  PIN f_mul_ex3_car[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 452.000 0.000 452.600 ;
    END
  END f_mul_ex3_car[2]
  PIN f_mul_ex3_car[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 456.000 0.000 456.600 ;
    END
  END f_mul_ex3_car[3]
  PIN f_mul_ex3_car[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 460.000 0.000 460.600 ;
    END
  END f_mul_ex3_car[4]
  PIN f_mul_ex3_car[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 464.000 0.000 464.600 ;
    END
  END f_mul_ex3_car[5]
  PIN f_mul_ex3_car[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 468.000 0.000 468.600 ;
    END
  END f_mul_ex3_car[6]
  PIN f_mul_ex3_car[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 472.000 0.000 472.600 ;
    END
  END f_mul_ex3_car[7]
  PIN f_mul_ex3_car[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 476.000 0.000 476.600 ;
    END
  END f_mul_ex3_car[8]
  PIN f_mul_ex3_car[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 480.000 0.000 480.600 ;
    END
  END f_mul_ex3_car[9]
  PIN f_mul_ex3_car[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 484.000 0.000 484.600 ;
    END
  END f_mul_ex3_car[10]
  PIN f_mul_ex3_car[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 488.000 0.000 488.600 ;
    END
  END f_mul_ex3_car[11]
  PIN f_mul_ex3_car[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 492.000 0.000 492.600 ;
    END
  END f_mul_ex3_car[12]
  PIN f_mul_ex3_car[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 496.000 0.000 496.600 ;
    END
  END f_mul_ex3_car[13]
  PIN f_mul_ex3_car[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 500.000 0.000 500.600 ;
    END
  END f_mul_ex3_car[14]
  PIN f_mul_ex3_car[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 504.000 0.000 504.600 ;
    END
  END f_mul_ex3_car[15]
  PIN f_mul_ex3_car[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 508.000 0.000 508.600 ;
    END
  END f_mul_ex3_car[16]
  PIN f_mul_ex3_car[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 512.000 0.000 512.600 ;
    END
  END f_mul_ex3_car[17]
  PIN f_mul_ex3_car[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 516.000 0.000 516.600 ;
    END
  END f_mul_ex3_car[18]
  PIN f_mul_ex3_car[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 520.000 0.000 520.600 ;
    END
  END f_mul_ex3_car[19]
  PIN f_mul_ex3_car[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 524.000 0.000 524.600 ;
    END
  END f_mul_ex3_car[20]
  PIN f_mul_ex3_car[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 528.000 0.000 528.600 ;
    END
  END f_mul_ex3_car[21]
  PIN f_mul_ex3_car[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 532.000 0.000 532.600 ;
    END
  END f_mul_ex3_car[22]
  PIN f_mul_ex3_car[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 536.000 0.000 536.600 ;
    END
  END f_mul_ex3_car[23]
  PIN f_mul_ex3_car[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 540.000 0.000 540.600 ;
    END
  END f_mul_ex3_car[24]
  PIN f_mul_ex3_car[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 544.000 0.000 544.600 ;
    END
  END f_mul_ex3_car[25]
  PIN f_mul_ex3_car[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 548.000 0.000 548.600 ;
    END
  END f_mul_ex3_car[26]
  PIN f_mul_ex3_car[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 552.000 0.000 552.600 ;
    END
  END f_mul_ex3_car[27]
  PIN f_mul_ex3_car[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 556.000 0.000 556.600 ;
    END
  END f_mul_ex3_car[28]
  PIN f_mul_ex3_car[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 560.000 0.000 560.600 ;
    END
  END f_mul_ex3_car[29]
  PIN f_mul_ex3_car[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 564.000 0.000 564.600 ;
    END
  END f_mul_ex3_car[30]
  PIN f_mul_ex3_car[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 568.000 0.000 568.600 ;
    END
  END f_mul_ex3_car[31]
  PIN f_mul_ex3_car[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 572.000 0.000 572.600 ;
    END
  END f_mul_ex3_car[32]
  PIN f_mul_ex3_car[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 576.000 0.000 576.600 ;
    END
  END f_mul_ex3_car[33]
  PIN f_mul_ex3_car[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 580.000 0.000 580.600 ;
    END
  END f_mul_ex3_car[34]
  PIN f_mul_ex3_car[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 584.000 0.000 584.600 ;
    END
  END f_mul_ex3_car[35]
  PIN f_mul_ex3_car[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 588.000 0.000 588.600 ;
    END
  END f_mul_ex3_car[36]
  PIN f_mul_ex3_car[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 592.000 0.000 592.600 ;
    END
  END f_mul_ex3_car[37]
  PIN f_mul_ex3_car[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 596.000 0.000 596.600 ;
    END
  END f_mul_ex3_car[38]
  PIN f_mul_ex3_car[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 600.000 0.000 600.600 ;
    END
  END f_mul_ex3_car[39]
  PIN f_mul_ex3_car[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 604.000 0.000 604.600 ;
    END
  END f_mul_ex3_car[40]
  PIN f_mul_ex3_car[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 608.000 0.000 608.600 ;
    END
  END f_mul_ex3_car[41]
  PIN f_mul_ex3_car[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 612.000 0.000 612.600 ;
    END
  END f_mul_ex3_car[42]
  PIN f_mul_ex3_car[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 616.000 0.000 616.600 ;
    END
  END f_mul_ex3_car[43]
  PIN f_mul_ex3_car[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 620.000 0.000 620.600 ;
    END
  END f_mul_ex3_car[44]
  PIN f_mul_ex3_car[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 624.000 0.000 624.600 ;
    END
  END f_mul_ex3_car[45]
  PIN f_mul_ex3_car[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 628.000 0.000 628.600 ;
    END
  END f_mul_ex3_car[46]
  PIN f_mul_ex3_car[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 632.000 0.000 632.600 ;
    END
  END f_mul_ex3_car[47]
  PIN f_mul_ex3_car[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 636.000 0.000 636.600 ;
    END
  END f_mul_ex3_car[48]
  PIN f_mul_ex3_car[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 640.000 0.000 640.600 ;
    END
  END f_mul_ex3_car[49]
  PIN f_mul_ex3_car[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 644.000 0.000 644.600 ;
    END
  END f_mul_ex3_car[50]
  PIN f_mul_ex3_car[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 648.000 0.000 648.600 ;
    END
  END f_mul_ex3_car[51]
  PIN f_mul_ex3_car[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 652.000 0.000 652.600 ;
    END
  END f_mul_ex3_car[52]
  PIN f_mul_ex3_car[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 656.000 0.000 656.600 ;
    END
  END f_mul_ex3_car[53]
  PIN f_mul_ex3_car[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 660.000 0.000 660.600 ;
    END
  END f_mul_ex3_car[54]
  PIN f_mul_ex3_car[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 664.000 0.000 664.600 ;
    END
  END f_mul_ex3_car[55]
  PIN f_mul_ex3_car[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 668.000 0.000 668.600 ;
    END
  END f_mul_ex3_car[56]
  PIN f_mul_ex3_car[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 672.000 0.000 672.600 ;
    END
  END f_mul_ex3_car[57]
  PIN f_mul_ex3_car[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 676.000 0.000 676.600 ;
    END
  END f_mul_ex3_car[58]
  PIN f_mul_ex3_car[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 680.000 0.000 680.600 ;
    END
  END f_mul_ex3_car[59]
  PIN f_mul_ex3_car[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 684.000 0.000 684.600 ;
    END
  END f_mul_ex3_car[60]
  PIN f_mul_ex3_car[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 688.000 0.000 688.600 ;
    END
  END f_mul_ex3_car[61]
  PIN f_mul_ex3_car[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 692.000 0.000 692.600 ;
    END
  END f_mul_ex3_car[62]
  PIN f_mul_ex3_car[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 696.000 0.000 696.600 ;
    END
  END f_mul_ex3_car[63]
  PIN f_mul_ex3_car[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 700.000 0.000 700.600 ;
    END
  END f_mul_ex3_car[64]
  PIN f_mul_ex3_car[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 704.000 0.000 704.600 ;
    END
  END f_mul_ex3_car[65]
  PIN f_mul_ex3_car[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 708.000 0.000 708.600 ;
    END
  END f_mul_ex3_car[66]
  PIN f_mul_ex3_car[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 712.000 0.000 712.600 ;
    END
  END f_mul_ex3_car[67]
  PIN f_mul_ex3_car[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 716.000 0.000 716.600 ;
    END
  END f_mul_ex3_car[68]
  PIN f_mul_ex3_car[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 720.000 0.000 720.600 ;
    END
  END f_mul_ex3_car[69]
  PIN f_mul_ex3_car[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 724.000 0.000 724.600 ;
    END
  END f_mul_ex3_car[70]
  PIN f_mul_ex3_car[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 728.000 0.000 728.600 ;
    END
  END f_mul_ex3_car[71]
  PIN f_mul_ex3_car[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 732.000 0.000 732.600 ;
    END
  END f_mul_ex3_car[72]
  PIN f_mul_ex3_car[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 736.000 0.000 736.600 ;
    END
  END f_mul_ex3_car[73]
  PIN f_mul_ex3_car[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 740.000 0.000 740.600 ;
    END
  END f_mul_ex3_car[74]
  PIN f_mul_ex3_car[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 744.000 0.000 744.600 ;
    END
  END f_mul_ex3_car[75]
  PIN f_mul_ex3_car[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 748.000 0.000 748.600 ;
    END
  END f_mul_ex3_car[76]
  PIN f_mul_ex3_car[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 752.000 0.000 752.600 ;
    END
  END f_mul_ex3_car[77]
  PIN f_mul_ex3_car[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 756.000 0.000 756.600 ;
    END
  END f_mul_ex3_car[78]
  PIN f_mul_ex3_car[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 760.000 0.000 760.600 ;
    END
  END f_mul_ex3_car[79]
  PIN f_mul_ex3_car[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 764.000 0.000 764.600 ;
    END
  END f_mul_ex3_car[80]
  PIN f_mul_ex3_car[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 768.000 0.000 768.600 ;
    END
  END f_mul_ex3_car[81]
  PIN f_mul_ex3_car[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 772.000 0.000 772.600 ;
    END
  END f_mul_ex3_car[82]
  PIN f_mul_ex3_car[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 776.000 0.000 776.600 ;
    END
  END f_mul_ex3_car[83]
  PIN f_mul_ex3_car[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 780.000 0.000 780.600 ;
    END
  END f_mul_ex3_car[84]
  PIN f_mul_ex3_car[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 784.000 0.000 784.600 ;
    END
  END f_mul_ex3_car[85]
  PIN f_mul_ex3_car[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 788.000 0.000 788.600 ;
    END
  END f_mul_ex3_car[86]
  PIN f_mul_ex3_car[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 792.000 0.000 792.600 ;
    END
  END f_mul_ex3_car[87]
  PIN f_mul_ex3_car[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 796.000 0.000 796.600 ;
    END
  END f_mul_ex3_car[88]
  PIN f_mul_ex3_car[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 800.000 0.000 800.600 ;
    END
  END f_mul_ex3_car[89]
  PIN f_mul_ex3_car[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 804.000 0.000 804.600 ;
    END
  END f_mul_ex3_car[90]
  PIN f_mul_ex3_car[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 808.000 0.000 808.600 ;
    END
  END f_mul_ex3_car[91]
  PIN f_mul_ex3_car[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 812.000 0.000 812.600 ;
    END
  END f_mul_ex3_car[92]
  PIN f_mul_ex3_car[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 816.000 0.000 816.600 ;
    END
  END f_mul_ex3_car[93]
  PIN f_mul_ex3_car[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 820.000 0.000 820.600 ;
    END
  END f_mul_ex3_car[94]
  PIN f_mul_ex3_car[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 824.000 0.000 824.600 ;
    END
  END f_mul_ex3_car[95]
  PIN f_mul_ex3_car[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 828.000 0.000 828.600 ;
    END
  END f_mul_ex3_car[96]
  PIN f_mul_ex3_car[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 832.000 0.000 832.600 ;
    END
  END f_mul_ex3_car[97]
  PIN f_mul_ex3_car[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 836.000 0.000 836.600 ;
    END
  END f_mul_ex3_car[98]
  PIN f_mul_ex3_car[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 840.000 0.000 840.600 ;
    END
  END f_mul_ex3_car[99]
  PIN f_mul_ex3_car[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 844.000 0.000 844.600 ;
    END
  END f_mul_ex3_car[100]
  PIN f_mul_ex3_car[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 848.000 0.000 848.600 ;
    END
  END f_mul_ex3_car[101]
  PIN f_mul_ex3_car[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 852.000 0.000 852.600 ;
    END
  END f_mul_ex3_car[102]
  PIN f_mul_ex3_car[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 856.000 0.000 856.600 ;
    END
  END f_mul_ex3_car[103]
  PIN f_mul_ex3_car[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 860.000 0.000 860.600 ;
    END
  END f_mul_ex3_car[104]
  PIN f_mul_ex3_car[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 864.000 0.000 864.600 ;
    END
  END f_mul_ex3_car[105]
  PIN f_mul_ex3_car[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 868.000 0.000 868.600 ;
    END
  END f_mul_ex3_car[106]
  PIN f_mul_ex3_car[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 872.000 0.000 872.600 ;
    END
  END f_mul_ex3_car[107]
  PIN f_mul_ex3_car[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.000 876.000 0.000 876.600 ;
    END
  END f_mul_ex3_car[108]
END tri_fu_mul
END LIBRARY

